module TOP #(parameter I=19, parameter F=11)
(
	input wire CLK,
	input wire RST, 
	input wire EN,
	
	input wire signed [I+F-1:0] IN0,
	input wire signed [I+F-1:0] IN1,
	input wire signed [I+F-1:0] IN2,
	input wire signed [I+F-1:0] IN3,
	input wire signed [I+F-1:0] IN4,
	input wire signed [I+F-1:0] IN5,
	input wire signed [I+F-1:0] IN6,
	input wire signed [I+F-1:0] IN7,
	input wire signed [I+F-1:0] IN8,
	input wire signed [I+F-1:0] IN9,
	input wire signed [I+F-1:0] IN10,
	input wire signed [I+F-1:0] IN11,
	input wire signed [I+F-1:0] IN12,
	input wire signed [I+F-1:0] IN13,
	input wire signed [I+F-1:0] IN14,
	input wire signed [I+F-1:0] IN15,
	input wire signed [I+F-1:0] IN16,
	input wire signed [I+F-1:0] IN17,
	input wire signed [I+F-1:0] IN18,
	input wire signed [I+F-1:0] IN19,
	input wire signed [I+F-1:0] IN20,
	input wire signed [I+F-1:0] IN21,
	input wire signed [I+F-1:0] IN22,
	input wire signed [I+F-1:0] IN23,
	input wire signed [I+F-1:0] IN24,
	input wire signed [I+F-1:0] IN25,
	input wire signed [I+F-1:0] IN26,
	input wire signed [I+F-1:0] IN27,
	input wire signed [I+F-1:0] IN28,
	input wire signed [I+F-1:0] IN29,
	input wire signed [I+F-1:0] IN30,
	input wire signed [I+F-1:0] IN31,
	
	output wire signed [I+F-1:0] OUT0_r,
	output wire signed [I+F-1:0] OUT0_i,
	output wire signed [I+F-1:0] OUT1_r,
	output wire signed [I+F-1:0] OUT1_i,
	output wire signed [I+F-1:0] OUT2_r,
	output wire signed [I+F-1:0] OUT2_i,
	output wire signed [I+F-1:0] OUT3_r,
	output wire signed [I+F-1:0] OUT3_i,
	output wire signed [I+F-1:0] OUT4_i,
	output wire signed [I+F-1:0] OUT4_r,
	output wire signed [I+F-1:0] OUT5_i,
	output wire signed [I+F-1:0] OUT5_r,
	output wire signed [I+F-1:0] OUT6_i,
	output wire signed [I+F-1:0] OUT6_r,
	output wire signed [I+F-1:0] OUT7_i,
	output wire signed [I+F-1:0] OUT7_r,
	output wire signed [I+F-1:0] OUT8_i,
	output wire signed [I+F-1:0] OUT8_r,
	output wire signed [I+F-1:0] OUT9_i,
	output wire signed [I+F-1:0] OUT9_r,
	output wire signed [I+F-1:0] OUT10_i,
	output wire signed [I+F-1:0] OUT10_r,
	output wire signed [I+F-1:0] OUT11_i,
	output wire signed [I+F-1:0] OUT11_r,
	output wire signed [I+F-1:0] OUT12_i,
	output wire signed [I+F-1:0] OUT12_r,
	output wire signed [I+F-1:0] OUT13_i,
	output wire signed [I+F-1:0] OUT13_r,
	output wire signed [I+F-1:0] OUT14_i,
	output wire signed [I+F-1:0] OUT14_r,
	output wire signed [I+F-1:0] OUT15_i,
	output wire signed [I+F-1:0] OUT15_r,
	output wire signed [I+F-1:0] OUT16_i,
	output wire signed [I+F-1:0] OUT16_r,
	output wire signed [I+F-1:0] OUT17_i,
	output wire signed [I+F-1:0] OUT17_r,
	output wire signed [I+F-1:0] OUT18_i,
	output wire signed [I+F-1:0] OUT18_r,
	output wire signed [I+F-1:0] OUT19_r,
	output wire signed [I+F-1:0] OUT19_i,
	output wire signed [I+F-1:0] OUT20_r,
	output wire signed [I+F-1:0] OUT20_i,
	output wire signed [I+F-1:0] OUT21_r,
	output wire signed [I+F-1:0] OUT21_i,
	output wire signed [I+F-1:0] OUT22_r,
	output wire signed [I+F-1:0] OUT22_i,
	output wire signed [I+F-1:0] OUT23_i,
	output wire signed [I+F-1:0] OUT23_r,
	output wire signed [I+F-1:0] OUT24_i,
	output wire signed [I+F-1:0] OUT24_r,
	output wire signed [I+F-1:0] OUT25_i,
	output wire signed [I+F-1:0] OUT25_r,
	output wire signed [I+F-1:0] OUT26_i,
	output wire signed [I+F-1:0] OUT26_r,
	output wire signed [I+F-1:0] OUT27_i,
	output wire signed [I+F-1:0] OUT27_r,
	output wire signed [I+F-1:0] OUT28_i,
	output wire signed [I+F-1:0] OUT28_r,
	output wire signed [I+F-1:0] OUT29_i,
	output wire signed [I+F-1:0] OUT29_r,
	output wire signed [I+F-1:0] OUT30_i,
	output wire signed [I+F-1:0] OUT30_r,
	output wire signed [I+F-1:0] OUT31_i,
	output wire signed [I+F-1:0] OUT31_r
	);
	


	reg signed [I+F-1:0] MAC0_IN1_R;
	reg signed [I+F-1:0] MAC0_IN1_I;
	reg signed [I+F-1:0] MAC0_IN2_R;
	reg signed [I+F-1:0] MAC0_IN2_I;
	reg signed [I+F-1:0] MAC1_IN1_R;
	reg signed [I+F-1:0] MAC1_IN1_I;
	reg signed [I+F-1:0] MAC1_IN2_R;
	reg signed [I+F-1:0] MAC1_IN2_I;
	reg signed [I+F-1:0] MAC2_IN1_R;
	reg signed [I+F-1:0] MAC2_IN1_I;
	reg signed [I+F-1:0] MAC2_IN2_R;
	reg signed [I+F-1:0] MAC2_IN2_I;
	reg signed [I+F-1:0] MAC3_IN1_R;
	reg signed [I+F-1:0] MAC3_IN1_I;
	reg signed [I+F-1:0] MAC3_IN2_R;
	reg signed [I+F-1:0] MAC3_IN2_I;
	reg signed [I+F-1:0] MAC4_IN1_R;
	reg signed [I+F-1:0] MAC4_IN1_I;
	reg signed [I+F-1:0] MAC4_IN2_R;
	reg signed [I+F-1:0] MAC4_IN2_I;
	reg signed [I+F-1:0] MAC5_IN1_R;
	reg signed [I+F-1:0] MAC5_IN1_I;
	reg signed [I+F-1:0] MAC5_IN2_R;
	reg signed [I+F-1:0] MAC5_IN2_I;
	reg signed [I+F-1:0] MAC6_IN1_R;
	reg signed [I+F-1:0] MAC6_IN1_I;
	reg signed [I+F-1:0] MAC6_IN2_R;
	reg signed [I+F-1:0] MAC6_IN2_I;
	reg signed [I+F-1:0] MAC7_IN1_R;
	reg signed [I+F-1:0] MAC7_IN1_I;
	reg signed [I+F-1:0] MAC7_IN2_R;
	reg signed [I+F-1:0] MAC7_IN2_I;
	reg signed [I+F-1:0] MAC8_IN1_R;
	reg signed [I+F-1:0] MAC8_IN1_I;
	reg signed [I+F-1:0] MAC8_IN2_R;
	reg signed [I+F-1:0] MAC8_IN2_I;
	reg signed [I+F-1:0] MAC9_IN1_R;
	reg signed [I+F-1:0] MAC9_IN1_I;
	reg signed [I+F-1:0] MAC9_IN2_R;
	reg signed [I+F-1:0] MAC9_IN2_I;
	reg signed [I+F-1:0] MAC10_IN1_R;
	reg signed [I+F-1:0] MAC10_IN1_I;
	reg signed [I+F-1:0] MAC10_IN2_R;
	reg signed [I+F-1:0] MAC10_IN2_I;
	reg signed [I+F-1:0] MAC11_IN1_R;
	reg signed [I+F-1:0] MAC11_IN1_I;
	reg signed [I+F-1:0] MAC11_IN2_R;
	reg signed [I+F-1:0] MAC11_IN2_I;
	reg signed [I+F-1:0] MAC12_IN1_R;
	reg signed [I+F-1:0] MAC12_IN1_I;
	reg signed [I+F-1:0] MAC12_IN2_R;
	reg signed [I+F-1:0] MAC12_IN2_I;
	reg signed [I+F-1:0] MAC13_IN1_R;
	reg signed [I+F-1:0] MAC13_IN1_I;
	reg signed [I+F-1:0] MAC13_IN2_R;
	reg signed [I+F-1:0] MAC13_IN2_I;
	reg signed [I+F-1:0] MAC14_IN1_R;
	reg signed [I+F-1:0] MAC14_IN1_I;
	reg signed [I+F-1:0] MAC14_IN2_R;
	reg signed [I+F-1:0] MAC14_IN2_I;
	reg signed [I+F-1:0] MAC15_IN1_R;
	reg signed [I+F-1:0] MAC15_IN1_I;
	reg signed [I+F-1:0] MAC15_IN2_R;
	reg signed [I+F-1:0] MAC15_IN2_I;



	wire signed [I+F-1:0] MAC0_OUT1_R;
	wire signed [I+F-1:0] MAC0_OUT1_I;
	wire signed [I+F-1:0] MAC0_OUT2_R;
	wire signed [I+F-1:0] MAC0_OUT2_I;
	wire signed [I+F-1:0] MAC1_OUT1_R;
	wire signed [I+F-1:0] MAC1_OUT1_I;
	wire signed [I+F-1:0] MAC1_OUT2_R;
	wire signed [I+F-1:0] MAC1_OUT2_I;
	wire signed [I+F-1:0] MAC2_OUT1_R;
	wire signed [I+F-1:0] MAC2_OUT1_I;
	wire signed [I+F-1:0] MAC2_OUT2_R;
	wire signed [I+F-1:0] MAC2_OUT2_I;
	wire signed [I+F-1:0] MAC3_OUT1_R;
	wire signed [I+F-1:0] MAC3_OUT1_I;
	wire signed [I+F-1:0] MAC3_OUT2_R;
	wire signed [I+F-1:0] MAC3_OUT2_I;
	wire signed [I+F-1:0] MAC4_OUT1_R;
	wire signed [I+F-1:0] MAC4_OUT1_I;
	wire signed [I+F-1:0] MAC4_OUT2_R;
	wire signed [I+F-1:0] MAC4_OUT2_I;
	wire signed [I+F-1:0] MAC5_OUT1_R;
	wire signed [I+F-1:0] MAC5_OUT1_I;
	wire signed [I+F-1:0] MAC5_OUT2_R;
	wire signed [I+F-1:0] MAC5_OUT2_I;
	wire signed [I+F-1:0] MAC6_OUT1_R;
	wire signed [I+F-1:0] MAC6_OUT1_I;
	wire signed [I+F-1:0] MAC6_OUT2_R;
	wire signed [I+F-1:0] MAC6_OUT2_I;
	wire signed [I+F-1:0] MAC7_OUT1_R;
	wire signed [I+F-1:0] MAC7_OUT1_I;
	wire signed [I+F-1:0] MAC7_OUT2_R;
	wire signed [I+F-1:0] MAC7_OUT2_I;
	wire signed [I+F-1:0] MAC8_OUT1_R;
	wire signed [I+F-1:0] MAC8_OUT1_I;
	wire signed [I+F-1:0] MAC8_OUT2_R;
	wire signed [I+F-1:0] MAC8_OUT2_I;
	wire signed [I+F-1:0] MAC9_OUT1_R;
	wire signed [I+F-1:0] MAC9_OUT1_I;
	wire signed [I+F-1:0] MAC9_OUT2_R;
	wire signed [I+F-1:0] MAC9_OUT2_I;
	wire signed [I+F-1:0] MAC10_OUT1_R;
	wire signed [I+F-1:0] MAC10_OUT1_I;
	wire signed [I+F-1:0] MAC10_OUT2_R;
	wire signed [I+F-1:0] MAC10_OUT2_I;
	wire signed [I+F-1:0] MAC11_OUT1_R;
	wire signed [I+F-1:0] MAC11_OUT1_I;
	wire signed [I+F-1:0] MAC11_OUT2_R;
	wire signed [I+F-1:0] MAC11_OUT2_I;
	wire signed [I+F-1:0] MAC12_OUT1_R;
	wire signed [I+F-1:0] MAC12_OUT1_I;
	wire signed [I+F-1:0] MAC12_OUT2_R;
	wire signed [I+F-1:0] MAC12_OUT2_I;
	wire signed [I+F-1:0] MAC13_OUT1_R;
	wire signed [I+F-1:0] MAC13_OUT1_I;
	wire signed [I+F-1:0] MAC13_OUT2_R;
	wire signed [I+F-1:0] MAC13_OUT2_I;
	wire signed [I+F-1:0] MAC14_OUT1_R;
	wire signed [I+F-1:0] MAC14_OUT1_I;
	wire signed [I+F-1:0] MAC14_OUT2_R;
	wire signed [I+F-1:0] MAC14_OUT2_I;
	wire signed [I+F-1:0] MAC15_OUT1_R;
	wire signed [I+F-1:0] MAC15_OUT1_I;
	wire signed [I+F-1:0] MAC15_OUT2_R;
	wire signed [I+F-1:0] MAC15_OUT2_I;
	
	reg signed [I+F-1:0] MAC0_W_R;
	reg signed [I+F-1:0] MAC0_W_I;
	reg signed [I+F-1:0] MAC1_W_R;
	reg signed [I+F-1:0] MAC1_W_I;
	reg signed [I+F-1:0] MAC2_W_R;
	reg signed [I+F-1:0] MAC2_W_I;
	reg signed [I+F-1:0] MAC3_W_R;
	reg signed [I+F-1:0] MAC3_W_I;
	reg signed [I+F-1:0] MAC4_W_R;
	reg signed [I+F-1:0] MAC4_W_I;
	reg signed [I+F-1:0] MAC5_W_R;
	reg signed [I+F-1:0] MAC5_W_I;
	reg signed [I+F-1:0] MAC6_W_R;
	reg signed [I+F-1:0] MAC6_W_I;
	reg signed [I+F-1:0] MAC7_W_R;
	reg signed [I+F-1:0] MAC7_W_I;
	reg signed [I+F-1:0] MAC8_W_R;
	reg signed [I+F-1:0] MAC8_W_I;
	reg signed [I+F-1:0] MAC9_W_R;
	reg signed [I+F-1:0] MAC9_W_I;
	reg signed [I+F-1:0] MAC10_W_R;
	reg signed [I+F-1:0] MAC10_W_I;
	reg signed [I+F-1:0] MAC11_W_R;
	reg signed [I+F-1:0] MAC11_W_I;
	reg signed [I+F-1:0] MAC12_W_R;
	reg signed [I+F-1:0] MAC12_W_I;
	reg signed [I+F-1:0] MAC13_W_R;
	reg signed [I+F-1:0] MAC13_W_I;
	reg signed [I+F-1:0] MAC14_W_R;
	reg signed [I+F-1:0] MAC14_W_I;
	reg signed [I+F-1:0] MAC15_W_R;
	reg signed [I+F-1:0] MAC15_W_I;
	
	
	wire signed [I+F-1:0] regfile0_out0_r;
	wire signed [I+F-1:0] regfile0_out0_i;
	wire signed [I+F-1:0] regfile0_out1_r;
	wire signed [I+F-1:0] regfile0_out1_i;
	wire signed [I+F-1:0] regfile0_out2_r;
	wire signed [I+F-1:0] regfile0_out2_i;
	wire signed [I+F-1:0] regfile0_out3_r;
	wire signed [I+F-1:0] regfile0_out3_i;
	wire signed [I+F-1:0] regfile0_out4_r;
	wire signed [I+F-1:0] regfile0_out4_i;
	wire signed [I+F-1:0] regfile0_out5_r;
	wire signed [I+F-1:0] regfile0_out5_i;
	wire signed [I+F-1:0] regfile0_out6_r;
	wire signed [I+F-1:0] regfile0_out6_i;
	wire signed [I+F-1:0] regfile0_out7_r;
	wire signed [I+F-1:0] regfile0_out7_i;
	wire signed [I+F-1:0] regfile0_out8_r;
	wire signed [I+F-1:0] regfile0_out8_i;
	wire signed [I+F-1:0] regfile0_out9_r;
	wire signed [I+F-1:0] regfile0_out9_i;
	wire signed [I+F-1:0] regfile0_out10_r;
	wire signed [I+F-1:0] regfile0_out10_i;
	wire signed [I+F-1:0] regfile0_out11_r;
	wire signed [I+F-1:0] regfile0_out11_i;
	wire signed [I+F-1:0] regfile0_out12_r;
	wire signed [I+F-1:0] regfile0_out12_i;
	wire signed [I+F-1:0] regfile0_out13_r;
	wire signed [I+F-1:0] regfile0_out13_i;
	wire signed [I+F-1:0] regfile0_out14_r;
	wire signed [I+F-1:0] regfile0_out14_i;
	wire signed [I+F-1:0] regfile0_out15_r;
	wire signed [I+F-1:0] regfile0_out15_i;
	wire signed [I+F-1:0] regfile0_out16_r;
	wire signed [I+F-1:0] regfile0_out16_i;
	wire signed [I+F-1:0] regfile0_out17_r;
	wire signed [I+F-1:0] regfile0_out17_i;
	wire signed [I+F-1:0] regfile0_out18_r;
	wire signed [I+F-1:0] regfile0_out18_i;
	wire signed [I+F-1:0] regfile0_out19_r;
	wire signed [I+F-1:0] regfile0_out19_i;
	wire signed [I+F-1:0] regfile0_out20_r;
	wire signed [I+F-1:0] regfile0_out20_i;
	wire signed [I+F-1:0] regfile0_out21_r;
	wire signed [I+F-1:0] regfile0_out21_i;
	wire signed [I+F-1:0] regfile0_out22_r;
	wire signed [I+F-1:0] regfile0_out22_i;
	wire signed [I+F-1:0] regfile0_out23_r;
	wire signed [I+F-1:0] regfile0_out23_i;
	wire signed [I+F-1:0] regfile0_out24_r;
	wire signed [I+F-1:0] regfile0_out24_i;
	wire signed [I+F-1:0] regfile0_out25_r;
	wire signed [I+F-1:0] regfile0_out25_i;
	wire signed [I+F-1:0] regfile0_out26_r;
	wire signed [I+F-1:0] regfile0_out26_i;
	wire signed [I+F-1:0] regfile0_out27_r;
	wire signed [I+F-1:0] regfile0_out27_i;
	wire signed [I+F-1:0] regfile0_out28_r;
	wire signed [I+F-1:0] regfile0_out28_i;
	wire signed [I+F-1:0] regfile0_out29_r;
	wire signed [I+F-1:0] regfile0_out29_i;
	wire signed [I+F-1:0] regfile0_out30_r;
	wire signed [I+F-1:0] regfile0_out30_i;
	wire signed [I+F-1:0] regfile0_out31_r;
	wire signed [I+F-1:0] regfile0_out31_i;
	
	wire signed [I+F-1:0] regfile1_out0_r;
	wire signed [I+F-1:0] regfile1_out0_i;
	wire signed [I+F-1:0] regfile1_out1_r;
	wire signed [I+F-1:0] regfile1_out1_i;
	wire signed [I+F-1:0] regfile1_out2_r;
	wire signed [I+F-1:0] regfile1_out2_i;
	wire signed [I+F-1:0] regfile1_out3_r;
	wire signed [I+F-1:0] regfile1_out3_i;
	wire signed [I+F-1:0] regfile1_out4_r;
	wire signed [I+F-1:0] regfile1_out4_i;
	wire signed [I+F-1:0] regfile1_out5_r;
	wire signed [I+F-1:0] regfile1_out5_i;
	wire signed [I+F-1:0] regfile1_out6_r;
	wire signed [I+F-1:0] regfile1_out6_i;
	wire signed [I+F-1:0] regfile1_out7_r;
	wire signed [I+F-1:0] regfile1_out7_i;
	wire signed [I+F-1:0] regfile1_out8_r;
	wire signed [I+F-1:0] regfile1_out8_i;
	wire signed [I+F-1:0] regfile1_out9_r;
	wire signed [I+F-1:0] regfile1_out9_i;
	wire signed [I+F-1:0] regfile1_out10_r;
	wire signed [I+F-1:0] regfile1_out10_i;
	wire signed [I+F-1:0] regfile1_out11_r;
	wire signed [I+F-1:0] regfile1_out11_i;
	wire signed [I+F-1:0] regfile1_out12_r;
	wire signed [I+F-1:0] regfile1_out12_i;
	wire signed [I+F-1:0] regfile1_out13_r;
	wire signed [I+F-1:0] regfile1_out13_i;
	wire signed [I+F-1:0] regfile1_out14_r;
	wire signed [I+F-1:0] regfile1_out14_i;
	wire signed [I+F-1:0] regfile1_out15_r;
	wire signed [I+F-1:0] regfile1_out15_i;
	wire signed [I+F-1:0] regfile1_out16_r;
	wire signed [I+F-1:0] regfile1_out16_i;
	wire signed [I+F-1:0] regfile1_out17_r;
	wire signed [I+F-1:0] regfile1_out17_i;
	wire signed [I+F-1:0] regfile1_out18_r;
	wire signed [I+F-1:0] regfile1_out18_i;
	wire signed [I+F-1:0] regfile1_out19_r;
	wire signed [I+F-1:0] regfile1_out19_i;
	wire signed [I+F-1:0] regfile1_out20_r;
	wire signed [I+F-1:0] regfile1_out20_i;
	wire signed [I+F-1:0] regfile1_out21_r;
	wire signed [I+F-1:0] regfile1_out21_i;
	wire signed [I+F-1:0] regfile1_out22_r;
	wire signed [I+F-1:0] regfile1_out22_i;
	wire signed [I+F-1:0] regfile1_out23_r;
	wire signed [I+F-1:0] regfile1_out23_i;
	wire signed [I+F-1:0] regfile1_out24_r;
	wire signed [I+F-1:0] regfile1_out24_i;
	wire signed [I+F-1:0] regfile1_out25_r;
	wire signed [I+F-1:0] regfile1_out25_i;
	wire signed [I+F-1:0] regfile1_out26_r;
	wire signed [I+F-1:0] regfile1_out26_i;
	wire signed [I+F-1:0] regfile1_out27_r;
	wire signed [I+F-1:0] regfile1_out27_i;
	wire signed [I+F-1:0] regfile1_out28_r;
	wire signed [I+F-1:0] regfile1_out28_i;
	wire signed [I+F-1:0] regfile1_out29_r;
	wire signed [I+F-1:0] regfile1_out29_i;
	wire signed [I+F-1:0] regfile1_out30_r;
	wire signed [I+F-1:0] regfile1_out30_i;
	wire signed [I+F-1:0] regfile1_out31_r;
	wire signed [I+F-1:0] regfile1_out31_i;
	
	wire signed [I+F-1:0] regfile2_out0_r;
	wire signed [I+F-1:0] regfile2_out0_i;
	wire signed [I+F-1:0] regfile2_out1_r;
	wire signed [I+F-1:0] regfile2_out1_i;
	wire signed [I+F-1:0] regfile2_out2_r;
	wire signed [I+F-1:0] regfile2_out2_i;
	wire signed [I+F-1:0] regfile2_out3_r;
	wire signed [I+F-1:0] regfile2_out3_i;
	wire signed [I+F-1:0] regfile2_out4_r;
	wire signed [I+F-1:0] regfile2_out4_i;
	wire signed [I+F-1:0] regfile2_out5_r;
	wire signed [I+F-1:0] regfile2_out5_i;
	wire signed [I+F-1:0] regfile2_out6_r;
	wire signed [I+F-1:0] regfile2_out6_i;
	wire signed [I+F-1:0] regfile2_out7_r;
	wire signed [I+F-1:0] regfile2_out7_i;
	wire signed [I+F-1:0] regfile2_out8_r;
	wire signed [I+F-1:0] regfile2_out8_i;
	wire signed [I+F-1:0] regfile2_out9_r;
	wire signed [I+F-1:0] regfile2_out9_i;
	wire signed [I+F-1:0] regfile2_out10_r;
	wire signed [I+F-1:0] regfile2_out10_i;
	wire signed [I+F-1:0] regfile2_out11_r;
	wire signed [I+F-1:0] regfile2_out11_i;
	wire signed [I+F-1:0] regfile2_out12_r;
	wire signed [I+F-1:0] regfile2_out12_i;
	wire signed [I+F-1:0] regfile2_out13_r;
	wire signed [I+F-1:0] regfile2_out13_i;
	wire signed [I+F-1:0] regfile2_out14_r;
	wire signed [I+F-1:0] regfile2_out14_i;
	wire signed [I+F-1:0] regfile2_out15_r;
	wire signed [I+F-1:0] regfile2_out15_i;
	wire signed [I+F-1:0] regfile2_out16_r;
	wire signed [I+F-1:0] regfile2_out16_i;
	wire signed [I+F-1:0] regfile2_out17_r;
	wire signed [I+F-1:0] regfile2_out17_i;
	wire signed [I+F-1:0] regfile2_out18_r;
	wire signed [I+F-1:0] regfile2_out18_i;
	wire signed [I+F-1:0] regfile2_out19_r;
	wire signed [I+F-1:0] regfile2_out19_i;
	wire signed [I+F-1:0] regfile2_out20_r;
	wire signed [I+F-1:0] regfile2_out20_i;
	wire signed [I+F-1:0] regfile2_out21_r;
	wire signed [I+F-1:0] regfile2_out21_i;
	wire signed [I+F-1:0] regfile2_out22_r;
	wire signed [I+F-1:0] regfile2_out22_i;
	wire signed [I+F-1:0] regfile2_out23_r;
	wire signed [I+F-1:0] regfile2_out23_i;
	wire signed [I+F-1:0] regfile2_out24_r;
	wire signed [I+F-1:0] regfile2_out24_i;
	wire signed [I+F-1:0] regfile2_out25_r;
	wire signed [I+F-1:0] regfile2_out25_i;
	wire signed [I+F-1:0] regfile2_out26_r;
	wire signed [I+F-1:0] regfile2_out26_i;
	wire signed [I+F-1:0] regfile2_out27_r;
	wire signed [I+F-1:0] regfile2_out27_i;
	wire signed [I+F-1:0] regfile2_out28_r;
	wire signed [I+F-1:0] regfile2_out28_i;
	wire signed [I+F-1:0] regfile2_out29_r;
	wire signed [I+F-1:0] regfile2_out29_i;
	wire signed [I+F-1:0] regfile2_out30_r;
	wire signed [I+F-1:0] regfile2_out30_i;
	wire signed [I+F-1:0] regfile2_out31_r;
	wire signed [I+F-1:0] regfile2_out31_i;
	
	wire signed [I+F-1:0] regfile3_out0_r;
	wire signed [I+F-1:0] regfile3_out0_i;
	wire signed [I+F-1:0] regfile3_out1_r;
	wire signed [I+F-1:0] regfile3_out1_i;
	wire signed [I+F-1:0] regfile3_out2_r;
	wire signed [I+F-1:0] regfile3_out2_i;
	wire signed [I+F-1:0] regfile3_out3_r;
	wire signed [I+F-1:0] regfile3_out3_i;
	wire signed [I+F-1:0] regfile3_out4_r;
	wire signed [I+F-1:0] regfile3_out4_i;
	wire signed [I+F-1:0] regfile3_out5_r;
	wire signed [I+F-1:0] regfile3_out5_i;
	wire signed [I+F-1:0] regfile3_out6_r;
	wire signed [I+F-1:0] regfile3_out6_i;
	wire signed [I+F-1:0] regfile3_out7_r;
	wire signed [I+F-1:0] regfile3_out7_i;
	wire signed [I+F-1:0] regfile3_out8_r;
	wire signed [I+F-1:0] regfile3_out8_i;
	wire signed [I+F-1:0] regfile3_out9_r;
	wire signed [I+F-1:0] regfile3_out9_i;
	wire signed [I+F-1:0] regfile3_out10_r;
	wire signed [I+F-1:0] regfile3_out10_i;
	wire signed [I+F-1:0] regfile3_out11_r;
	wire signed [I+F-1:0] regfile3_out11_i;
	wire signed [I+F-1:0] regfile3_out12_r;
	wire signed [I+F-1:0] regfile3_out12_i;
	wire signed [I+F-1:0] regfile3_out13_r;
	wire signed [I+F-1:0] regfile3_out13_i;
	wire signed [I+F-1:0] regfile3_out14_r;
	wire signed [I+F-1:0] regfile3_out14_i;
	wire signed [I+F-1:0] regfile3_out15_r;
	wire signed [I+F-1:0] regfile3_out15_i;
	wire signed [I+F-1:0] regfile3_out16_r;
	wire signed [I+F-1:0] regfile3_out16_i;
	wire signed [I+F-1:0] regfile3_out17_r;
	wire signed [I+F-1:0] regfile3_out17_i;
	wire signed [I+F-1:0] regfile3_out18_r;
	wire signed [I+F-1:0] regfile3_out18_i;
	wire signed [I+F-1:0] regfile3_out19_r;
	wire signed [I+F-1:0] regfile3_out19_i;
	wire signed [I+F-1:0] regfile3_out20_r;
	wire signed [I+F-1:0] regfile3_out20_i;
	wire signed [I+F-1:0] regfile3_out21_r;
	wire signed [I+F-1:0] regfile3_out21_i;
	wire signed [I+F-1:0] regfile3_out22_r;
	wire signed [I+F-1:0] regfile3_out22_i;
	wire signed [I+F-1:0] regfile3_out23_r;
	wire signed [I+F-1:0] regfile3_out23_i;
	wire signed [I+F-1:0] regfile3_out24_r;
	wire signed [I+F-1:0] regfile3_out24_i;
	wire signed [I+F-1:0] regfile3_out25_r;
	wire signed [I+F-1:0] regfile3_out25_i;
	wire signed [I+F-1:0] regfile3_out26_r;
	wire signed [I+F-1:0] regfile3_out26_i;
	wire signed [I+F-1:0] regfile3_out27_r;
	wire signed [I+F-1:0] regfile3_out27_i;
	wire signed [I+F-1:0] regfile3_out28_r;
	wire signed [I+F-1:0] regfile3_out28_i;
	wire signed [I+F-1:0] regfile3_out29_r;
	wire signed [I+F-1:0] regfile3_out29_i;
	wire signed [I+F-1:0] regfile3_out30_r;
	wire signed [I+F-1:0] regfile3_out30_i;
	wire signed [I+F-1:0] regfile3_out31_r;
	wire signed [I+F-1:0] regfile3_out31_i;
	
	wire  E0;
	wire  E1;
	wire  E2;
	wire  E3;
	wire  E4;
	
	wire [3:0] Sel;
	
always@(*)
begin
			if ( Sel == 4'd1)
				begin
						 MAC0_IN1_R<=IN0;
						 MAC0_IN1_I<=0;
						 MAC0_IN2_R<=IN16;
						 MAC0_IN2_I<=0;
						 MAC1_IN1_R<=IN8;
						 MAC1_IN1_I<=0;
						 MAC1_IN2_R<=IN24;
						 MAC1_IN2_I<=0;
						 MAC2_IN1_R<=IN4;
						 MAC2_IN1_I<=0;
						 MAC2_IN2_R<=IN20;
						 MAC2_IN2_I<=0;
						 MAC3_IN1_R<=IN12;
						 MAC3_IN1_I<=0;
						 MAC3_IN2_R<=IN28;
						 MAC3_IN2_I<=0;
						 MAC4_IN1_R<=IN2;
						 MAC4_IN1_I<=0;
						 MAC4_IN2_R<=IN14;
						 MAC4_IN2_I<=0;
						 MAC5_IN1_R<=IN10;
						 MAC5_IN1_I<=0;
						 MAC5_IN2_R<=IN26;
						 MAC5_IN2_I<=0;
						 MAC6_IN1_R<=IN6;
						 MAC6_IN1_I<=0;
						 MAC6_IN2_R<=IN22;
						 MAC6_IN2_I<=0;
						 MAC7_IN1_R<=IN14;
						 MAC7_IN1_I<=0;
						 MAC7_IN2_R<=IN30;
						 MAC7_IN2_I<=0;
						 MAC8_IN1_R<=IN1;
						 MAC8_IN1_I<=0;
						 MAC8_IN2_R<=IN17;
						 MAC8_IN2_I<=0;
						 MAC9_IN1_R<=IN9;
						 MAC9_IN1_I<=0;
						 MAC9_IN2_R<=IN25;
						 MAC9_IN2_I<=0;
						 MAC10_IN1_R<=IN5;
						 MAC10_IN1_I<=0;
						 MAC10_IN2_R<=IN21;
						 MAC10_IN2_I<=0;
						 MAC11_IN1_R<=IN13;
						 MAC11_IN1_I<=0;
						 MAC11_IN2_R<=IN29;
						 MAC11_IN2_I<=0;
						 MAC12_IN1_R<=IN3;
						 MAC12_IN1_I<=0;
						 MAC12_IN2_R<=IN19;
						 MAC12_IN2_I<=0;
						 MAC13_IN1_R<=IN11;
						 MAC13_IN1_I<=0;
						 MAC13_IN2_R<=IN27;
						 MAC13_IN2_I<=0;
						 MAC14_IN1_R<=IN7;
						 MAC14_IN1_I<=0;
						 MAC14_IN2_R<=IN23;
						 MAC14_IN2_I<=0;
						 MAC15_IN1_R<=IN15;
						 MAC15_IN1_I<=0;
						 MAC15_IN2_R<=IN31;
						 MAC15_IN2_I<=0;
						 
						 MAC0_W_R<=30'b000000000000000000100000000000;
						 MAC0_W_I<=0;
						 MAC1_W_R<=30'b000000000000000000100000000000;
						 MAC1_W_I<=0;
						 MAC2_W_R<=30'b000000000000000000100000000000;
						 MAC2_W_I<=0;
						 MAC3_W_R<=30'b000000000000000000100000000000;
						 MAC3_W_I<=0;
						 MAC4_W_R<=30'b000000000000000000100000000000;
						 MAC4_W_I<=0;
						 MAC5_W_R<=30'b000000000000000000100000000000;
						 MAC5_W_I<=0;
						 MAC6_W_R<=30'b000000000000000000100000000000;
						 MAC6_W_I<=0;
						 MAC7_W_R<=30'b000000000000000000100000000000;
						 MAC7_W_I<=0;
						 MAC8_W_R<=30'b000000000000000000100000000000;
						 MAC8_W_I<=0;
						 MAC9_W_R<=30'b000000000000000000100000000000;
						 MAC9_W_I<=0;
						 MAC10_W_R<=30'b000000000000000000100000000000;
						 MAC10_W_I<=0;
						 MAC11_W_R<=30'b000000000000000000100000000000;
						 MAC11_W_I<=0;
						 MAC12_W_R<=30'b000000000000000000100000000000;
						 MAC12_W_I<=0;
						 MAC13_W_R<=30'b000000000000000000100000000000;
						 MAC13_W_I<=0;
						 MAC14_W_R<=30'b000000000000000000100000000000;
						 MAC14_W_I<=0;
						 MAC15_W_R<=30'b000000000000000000100000000000;
						 MAC15_W_I<=0;		
				end
			else if	( Sel == 4'd2)
				begin
						 MAC0_IN1_R<=regfile0_out0_r;
						 MAC0_IN1_I<=regfile0_out0_i;
						 MAC0_IN2_R<=regfile0_out2_r;
						 MAC0_IN2_I<=regfile0_out2_i;
						 MAC1_IN1_R<=regfile0_out1_r;
						 MAC1_IN1_I<=regfile0_out1_i;
						 MAC1_IN2_R<=regfile0_out3_r;
						 MAC1_IN2_I<=regfile0_out3_i;
						 MAC2_IN1_R<=regfile0_out4_r;
						 MAC2_IN1_I<=regfile0_out4_i;
						 MAC2_IN2_R<=regfile0_out6_r;
						 MAC2_IN2_I<=regfile0_out6_i;
						 MAC3_IN1_R<=regfile0_out5_r;
						 MAC3_IN1_I<=regfile0_out5_i;
						 MAC3_IN2_R<=regfile0_out7_r;
						 MAC3_IN2_I<=regfile0_out7_i;
						 MAC4_IN1_R<=regfile0_out8_r;
						 MAC4_IN1_I<=regfile0_out8_i;
						 MAC4_IN2_R<=regfile0_out10_r;
						 MAC4_IN2_I<=regfile0_out10_i;
						 MAC5_IN1_R<=regfile0_out9_r;
						 MAC5_IN1_I<=regfile0_out9_i;
						 MAC5_IN2_R<=regfile0_out11_r;
						 MAC5_IN2_I<=regfile0_out11_i;
						 MAC6_IN1_R<=regfile0_out12_r;
						 MAC6_IN1_I<=regfile0_out12_i;
						 MAC6_IN2_R<=regfile0_out14_r;
						 MAC6_IN2_I<=regfile0_out14_i;
						 MAC7_IN1_R<=regfile0_out13_r;
						 MAC7_IN1_I<=regfile0_out13_i;
						 MAC7_IN2_R<=regfile0_out15_r;
						 MAC7_IN2_I<=regfile0_out15_i;
						 MAC8_IN1_R<=regfile0_out16_r;
						 MAC8_IN1_I<=regfile0_out16_i;
						 MAC8_IN2_R<=regfile0_out18_r;
						 MAC8_IN2_I<=regfile0_out18_i;
						 MAC9_IN1_R<=regfile0_out17_r;
						 MAC9_IN1_I<=regfile0_out17_i;
						 MAC9_IN2_R<=regfile0_out19_r;
						 MAC9_IN2_I<=regfile0_out19_i;
						 MAC10_IN1_R<=regfile0_out20_r;
						 MAC10_IN1_I<=regfile0_out20_i;
						 MAC10_IN2_R<=regfile0_out22_r;
						 MAC10_IN2_I<=regfile0_out22_i;
						 MAC11_IN1_R<=regfile0_out21_r;
						 MAC11_IN1_I<=regfile0_out21_i;
						 MAC11_IN2_R<=regfile0_out23_r;
						 MAC11_IN2_I<=regfile0_out23_i;
						 MAC12_IN1_R<=regfile0_out24_r;
						 MAC12_IN1_I<=regfile0_out24_i;
						 MAC12_IN2_R<=regfile0_out26_r;
						 MAC12_IN2_I<=regfile0_out26_i;
						 MAC13_IN1_R<=regfile0_out25_r;
						 MAC13_IN1_I<=regfile0_out25_i;
						 MAC13_IN2_R<=regfile0_out27_r;
						 MAC13_IN2_I<=regfile0_out27_i;
						 MAC14_IN1_R<=regfile0_out28_r;
						 MAC14_IN1_I<=regfile0_out28_i;
						 MAC14_IN2_R<=regfile0_out30_r;
						 MAC14_IN2_I<=regfile0_out30_i;
						 MAC15_IN1_R<=regfile0_out29_r;
						 MAC15_IN1_I<=regfile0_out29_i;
						 MAC15_IN2_R<=regfile0_out31_r;
						 MAC15_IN2_I<=regfile0_out31_i;
						 
						 MAC0_W_R<=30'b000000000000000000100000000000;
						 MAC0_W_I<=0;
						 MAC1_W_R<=0;
						 MAC1_W_I<=30'b111111111111111111100000000000;
						 MAC2_W_R<=30'b000000000000000000100000000000;
						 MAC2_W_I<=0;
						 MAC3_W_R<=0;
						 MAC3_W_I<=30'b111111111111111111100000000000;
						 MAC4_W_R<=30'b000000000000000000100000000000;
						 MAC4_W_I<=0;
						 MAC5_W_R<=0;
						 MAC5_W_I<=30'b111111111111111111100000000000;
						 MAC6_W_R<=30'b000000000000000000100000000000;
						 MAC6_W_I<=0;
						 MAC7_W_R<=0;
						 MAC7_W_I<=30'b111111111111111111100000000000;
						 MAC8_W_R<=30'b000000000000000000100000000000;
						 MAC8_W_I<=0;
						 MAC9_W_R<=0;
						 MAC9_W_I<=30'b111111111111111111100000000000;
						 MAC10_W_R<=30'b000000000000000000100000000000;
						 MAC10_W_I<=0;
						 MAC11_W_R<=0;
						 MAC11_W_I<=30'b111111111111111111100000000000;
						 MAC12_W_R<=30'b000000000000000000100000000000;
						 MAC12_W_I<=0;
						 MAC13_W_R<=0;
						 MAC13_W_I<=30'b111111111111111111100000000000;
						 MAC14_W_R<=30'b000000000000000000100000000000;
						 MAC14_W_I<=0;
						 MAC15_W_R<=0;
						 MAC15_W_I<=30'b111111111111111111100000000000;				
				end
			else if	( Sel == 4'd3)
				begin
						 MAC0_IN1_R<=regfile1_out0_r;
						 MAC0_IN1_I<=regfile1_out0_i;
						 MAC0_IN2_R<=regfile1_out4_r;
						 MAC0_IN2_I<=regfile1_out4_i;
						 MAC1_IN1_R<=regfile1_out1_r;
						 MAC1_IN1_I<=regfile1_out1_i;
						 MAC1_IN2_R<=regfile1_out5_r;
						 MAC1_IN2_I<=regfile1_out5_i;
						 MAC2_IN1_R<=regfile1_out2_r;
						 MAC2_IN1_I<=regfile1_out2_i;
						 MAC2_IN2_R<=regfile1_out6_r;
						 MAC2_IN2_I<=regfile1_out6_i;
						 MAC3_IN1_R<=regfile1_out3_r;
						 MAC3_IN1_I<=regfile1_out3_i;
						 MAC3_IN2_R<=regfile1_out7_r;
						 MAC3_IN2_I<=regfile1_out7_i;
						 MAC4_IN1_R<=regfile1_out8_r;
						 MAC4_IN1_I<=regfile1_out8_i;
						 MAC4_IN2_R<=regfile1_out12_r;
						 MAC4_IN2_I<=regfile1_out12_i;
						 MAC5_IN1_R<=regfile1_out9_r;
						 MAC5_IN1_I<=regfile1_out9_i;
						 MAC5_IN2_R<=regfile1_out13_r;
						 MAC5_IN2_I<=regfile1_out13_i;
						 MAC6_IN1_R<=regfile1_out10_r;
						 MAC6_IN1_I<=regfile1_out10_i;
						 MAC6_IN2_R<=regfile1_out14_r;
						 MAC6_IN2_I<=regfile1_out14_i;
						 MAC7_IN1_R<=regfile1_out11_r;
						 MAC7_IN1_I<=regfile1_out11_i;
						 MAC7_IN2_R<=regfile1_out15_r;
						 MAC7_IN2_I<=regfile1_out15_i;
						 MAC8_IN1_R<=regfile1_out16_r;
						 MAC8_IN1_I<=regfile1_out16_i;
						 MAC8_IN2_R<=regfile1_out20_r;
						 MAC8_IN2_I<=regfile1_out20_i;
						 MAC9_IN1_R<=regfile1_out17_r;
						 MAC9_IN1_I<=regfile1_out17_i;
						 MAC9_IN2_R<=regfile1_out21_r;
						 MAC9_IN2_I<=regfile1_out21_i;
						 MAC10_IN1_R<=regfile1_out18_r;
						 MAC10_IN1_I<=regfile1_out18_i;
						 MAC10_IN2_R<=regfile1_out22_r;
						 MAC10_IN2_I<=regfile1_out22_i;
						 MAC11_IN1_R<=regfile1_out19_r;
						 MAC11_IN1_I<=regfile1_out19_i;
						 MAC11_IN2_R<=regfile1_out23_r;
						 MAC11_IN2_I<=regfile1_out23_i;
						 MAC12_IN1_R<=regfile1_out24_r;
						 MAC12_IN1_I<=regfile1_out24_i;
						 MAC12_IN2_R<=regfile1_out28_r;
						 MAC12_IN2_I<=regfile1_out28_i;
						 MAC13_IN1_R<=regfile1_out25_r;
						 MAC13_IN1_I<=regfile1_out25_i;
						 MAC13_IN2_R<=regfile1_out29_r;
						 MAC13_IN2_I<=regfile1_out29_i;
						 MAC14_IN1_R<=regfile1_out26_r;
						 MAC14_IN1_I<=regfile1_out26_i;
						 MAC14_IN2_R<=regfile1_out30_r;
						 MAC14_IN2_I<=regfile1_out30_i;
						 MAC15_IN1_R<=regfile1_out27_r;
						 MAC15_IN1_I<=regfile1_out27_i;
						 MAC15_IN2_R<=regfile1_out31_r;
						 MAC15_IN2_I<=regfile1_out31_i;
						 
						 MAC0_W_R<=30'b000000000000000000100000000000;	
						 MAC0_W_I<=0;
						 MAC1_W_R<=30'b000000000000000000010110101000;
						 MAC1_W_I<=30'b111111111111111111101001011000;
						 MAC2_W_R<=0;
						 MAC2_W_I<=30'b111111111111111111100000000000;
						 MAC3_W_R<=30'b111111111111111111101001011000;
						 MAC3_W_I<=30'b111111111111111111101001011000;
						 MAC4_W_R<=30'b000000000000000000100000000000;	
						 MAC4_W_I<=0;
						 MAC5_W_R<=30'b000000000000000000010110101000;
						 MAC5_W_I<=30'b111111111111111111101001011000;
						 MAC6_W_R<=0;
						 MAC6_W_I<=30'b111111111111111111100000000000;
						 MAC7_W_R<=30'b111111111111111111101001011000;
						 MAC7_W_I<=30'b111111111111111111101001011000;
						 MAC8_W_R<=30'b000000000000000000100000000000;	
						 MAC8_W_I<=0;
						 MAC9_W_R<=30'b000000000000000000010110101000;
						 MAC9_W_I<=30'b111111111111111111101001011000;
						 MAC10_W_R<=0;
						 MAC10_W_I<=30'b111111111111111111100000000000;
						 MAC11_W_R<=30'b111111111111111111101001011000;
						 MAC11_W_I<=30'b111111111111111111101001011000;
						 MAC12_W_R<=30'b000000000000000000100000000000;	
						 MAC12_W_I<=0;
						 MAC13_W_R<=30'b000000000000000000010110101000;
						 MAC13_W_I<=30'b111111111111111111101001011000;
						 MAC14_W_R<=0;
						 MAC14_W_I<=30'b111111111111111111100000000000;
						 MAC15_W_R<=30'b111111111111111111101001011000;
						 MAC15_W_I<=30'b111111111111111111101001011000;		
				end
			else if	( Sel == 4'd4)
				begin
						MAC0_IN1_R<=regfile2_out0_r;
						 MAC0_IN1_I<=regfile2_out0_i;
						 MAC0_IN2_R<=regfile2_out8_r;
						 MAC0_IN2_I<=regfile2_out8_i;
						 MAC1_IN1_R<=regfile2_out1_r;
						 MAC1_IN1_I<=regfile2_out1_i;
						 MAC1_IN2_R<=regfile2_out9_r;
						 MAC1_IN2_I<=regfile2_out9_i;
						 MAC2_IN1_R<=regfile2_out2_r;
						 MAC2_IN1_I<=regfile2_out2_i;
						 MAC2_IN2_R<=regfile2_out10_r;
						 MAC2_IN2_I<=regfile2_out10_i;
						 MAC3_IN1_R<=regfile2_out3_r;
						 MAC3_IN1_I<=regfile2_out3_i;
						 MAC3_IN2_R<=regfile2_out11_r;
						 MAC3_IN2_I<=regfile2_out11_i;
						 MAC4_IN1_R<=regfile2_out4_r;
						 MAC4_IN1_I<=regfile2_out4_i;
						 MAC4_IN2_R<=regfile2_out12_r;
						 MAC4_IN2_I<=regfile2_out12_i;
						 MAC5_IN1_R<=regfile2_out5_r;
						 MAC5_IN1_I<=regfile2_out5_i;
						 MAC5_IN2_R<=regfile2_out13_r;
						 MAC5_IN2_I<=regfile2_out13_i;
						 MAC6_IN1_R<=regfile2_out6_r;
						 MAC6_IN1_I<=regfile2_out6_i;
						 MAC6_IN2_R<=regfile2_out14_r;
						 MAC6_IN2_I<=regfile2_out14_i;
						 MAC7_IN1_R<=regfile2_out7_r;
						 MAC7_IN1_I<=regfile2_out7_i;
						 MAC7_IN2_R<=regfile2_out15_r;
						 MAC7_IN2_I<=regfile2_out15_i;
						 MAC8_IN1_R<=regfile2_out16_r;
						 MAC8_IN1_I<=regfile2_out16_i;
						 MAC8_IN2_R<=regfile2_out24_r;
						 MAC8_IN2_I<=regfile2_out24_i;
						 MAC9_IN1_R<=regfile2_out17_r;
						 MAC9_IN1_I<=regfile2_out17_i;
						 MAC9_IN2_R<=regfile2_out25_r;
						 MAC9_IN2_I<=regfile2_out25_i;
						 MAC10_IN1_R<=regfile2_out18_r;
						 MAC10_IN1_I<=regfile2_out18_i;
						 MAC10_IN2_R<=regfile2_out26_r;
						 MAC10_IN2_I<=regfile2_out26_i;
						 MAC11_IN1_R<=regfile2_out19_r;
						 MAC11_IN1_I<=regfile2_out19_i;
						 MAC11_IN2_R<=regfile2_out27_r;
						 MAC11_IN2_I<=regfile2_out27_i;
						 MAC12_IN1_R<=regfile2_out20_r;
						 MAC12_IN1_I<=regfile2_out20_i;
						 MAC12_IN2_R<=regfile2_out28_r;
						 MAC12_IN2_I<=regfile2_out28_i;
						 MAC13_IN1_R<=regfile2_out21_r;
						 MAC13_IN1_I<=regfile2_out21_i;
						 MAC13_IN2_R<=regfile2_out29_r;
						 MAC13_IN2_I<=regfile2_out29_i;
						 MAC14_IN1_R<=regfile2_out22_r;
						 MAC14_IN1_I<=regfile2_out22_i;
						 MAC14_IN2_R<=regfile2_out30_r;
						 MAC14_IN2_I<=regfile2_out30_i;
						 MAC15_IN1_R<=regfile2_out23_r;
						 MAC15_IN1_I<=regfile2_out23_i;
						 MAC15_IN2_R<=regfile2_out31_r;
						 MAC15_IN2_I<=regfile2_out31_i;
						 
						 MAC0_W_R<=30'b000000000000000000100000000000;
						 MAC0_W_I<=0;
						 MAC1_W_R<=30'b000000000000000000011101100100;
						 MAC1_W_I<=30'b111111111111111111110011110000;
						 MAC2_W_R<=30'b000000000000000000010110101000;
						 MAC2_W_I<=30'b111111111111111111101001011000;
						 MAC3_W_R<=30'b000000000000000000001100010000;
						 MAC3_W_I<=30'b111111111111111111100010011100;
						 MAC4_W_R<=0;
						 MAC4_W_I<=30'b111111111111111111100000000000;
						 MAC5_W_R<=30'b111111111111111111110011110000;
						 MAC5_W_I<=30'b111111111111111111100010011100;
						 MAC6_W_R<=30'b111111111111111111101001011000;
						 MAC6_W_I<=30'b111111111111111111101001011000;
						 MAC7_W_R<=30'b111111111111111111100010011100;
						 MAC7_W_I<=30'b111111111111111111110011110000;
						 MAC8_W_R<=30'b000000000000000000100000000000;
						 MAC8_W_I<=0;
						 MAC9_W_R<=30'b000000000000000000011101100100;
						 MAC9_W_I<=30'b111111111111111111110011110000;
						 MAC10_W_R<=30'b000000000000000000010110101000;
						 MAC10_W_I<=30'b111111111111111111101001011000;
						 MAC11_W_R<=30'b000000000000000000001100010000;
						 MAC11_W_I<=30'b111111111111111111100010011100;
						 MAC12_W_R<=0;
						 MAC12_W_I<=30'b111111111111111111100000000000;
						 MAC13_W_R<=30'b111111111111111111110011110000;
						 MAC13_W_I<=30'b111111111111111111100010011100;
						 MAC14_W_R<=30'b111111111111111111101001011000;
						 MAC14_W_I<=30'b111111111111111111101001011000;
						 MAC15_W_R<=30'b111111111111111111100010011100;
						 MAC15_W_I<=30'b111111111111111111110011110000;
				end
			else if	( Sel == 4'd5)
				begin
						 MAC0_IN1_R<=regfile3_out0_r;
						 MAC0_IN1_I<=regfile3_out0_i;
						 MAC0_IN2_R<=regfile3_out8_r;
						 MAC0_IN2_I<=regfile3_out8_i;
						 MAC1_IN1_R<=regfile3_out1_r;
						 MAC1_IN1_I<=regfile3_out1_i;
						 MAC1_IN2_R<=regfile3_out9_r;
						 MAC1_IN2_I<=regfile3_out9_i;
						 MAC2_IN1_R<=regfile3_out2_r;
						 MAC2_IN1_I<=regfile3_out2_i;
						 MAC2_IN2_R<=regfile3_out10_r;
						 MAC2_IN2_I<=regfile3_out10_i;
						 MAC3_IN1_R<=regfile3_out3_r;
						 MAC3_IN1_I<=regfile3_out3_i;
						 MAC3_IN2_R<=regfile3_out11_r;
						 MAC3_IN2_I<=regfile3_out11_i;
						 MAC4_IN1_R<=regfile3_out4_r;
						 MAC4_IN1_I<=regfile3_out4_i;
						 MAC4_IN2_R<=regfile3_out12_r;
						 MAC4_IN2_I<=regfile3_out12_i;
						 MAC5_IN1_R<=regfile3_out5_r;
						 MAC5_IN1_I<=regfile3_out5_i;
						 MAC5_IN2_R<=regfile3_out13_r;
						 MAC5_IN2_I<=regfile3_out13_i;
						 MAC6_IN1_R<=regfile3_out6_r;
						 MAC6_IN1_I<=regfile3_out6_i;
						 MAC6_IN2_R<=regfile3_out14_r;
						 MAC6_IN2_I<=regfile3_out14_i;
						 MAC7_IN1_R<=regfile3_out7_r;
						 MAC7_IN1_I<=regfile3_out7_i;
						 MAC7_IN2_R<=regfile3_out15_r;
						 MAC7_IN2_I<=regfile3_out15_i;
						 MAC8_IN1_R<=regfile3_out16_r;
						 MAC8_IN1_I<=regfile3_out16_i;
						 MAC8_IN2_R<=regfile3_out24_r;
						 MAC8_IN2_I<=regfile3_out24_i;
						 MAC9_IN1_R<=regfile3_out17_r;
						 MAC9_IN1_I<=regfile3_out17_i;
						 MAC9_IN2_R<=regfile3_out25_r;
						 MAC9_IN2_I<=regfile3_out25_i;
						 MAC10_IN1_R<=regfile3_out18_r;
						 MAC10_IN1_I<=regfile3_out18_i;
						 MAC10_IN2_R<=regfile3_out26_r;
						 MAC10_IN2_I<=regfile3_out26_i;
						 MAC11_IN1_R<=regfile3_out19_r;
						 MAC11_IN1_I<=regfile3_out19_i;
						 MAC11_IN2_R<=regfile3_out27_r;
						 MAC11_IN2_I<=regfile3_out27_i;
						 MAC12_IN1_R<=regfile3_out20_r;
						 MAC12_IN1_I<=regfile3_out20_i;
						 MAC12_IN2_R<=regfile3_out28_r;
						 MAC12_IN2_I<=regfile3_out28_i;
						 MAC13_IN1_R<=regfile3_out21_r;
						 MAC13_IN1_I<=regfile3_out21_i;
						 MAC13_IN2_R<=regfile3_out29_r;
						 MAC13_IN2_I<=regfile3_out29_i;
						 MAC14_IN1_R<=regfile3_out22_r;
						 MAC14_IN1_I<=regfile3_out22_i;
						 MAC14_IN2_R<=regfile3_out30_r;
						 MAC14_IN2_I<=regfile3_out30_i;
						 MAC15_IN1_R<=regfile3_out23_r;
						 MAC15_IN1_I<=regfile3_out23_i;
						 MAC15_IN2_R<=regfile3_out31_r;
						 MAC15_IN2_I<=regfile3_out31_i;
						 
						 MAC0_W_R<=30'b000000000000000000100000000000;
						 MAC0_W_I<=0;
						 MAC1_W_R<=30'b000000000000000000011111011001;
						 MAC1_W_I<=30'b111111111111111111111001110000;
						 MAC2_W_R<=30'b000000000000000000011101100100;
						 MAC2_W_I<=30'b111111111111111111110011110000;
						 MAC3_W_R<=30'b000000000000000000011010100111;
						 MAC3_W_I<=30'b111111111111111111101110001110;
						 MAC4_W_R<=30'b000000000000000000010110101000;
						 MAC4_W_I<=30'b111111111111111111101001011000;
						 MAC5_W_R<=30'b000000000000000000010001110010;
						 MAC5_W_I<=30'b111111111111111111100101011001;
						 MAC6_W_R<=30'b000000000000000000001100010000;
						 MAC6_W_I<=30'b111111111111111111100010011100;
						 MAC7_W_R<=30'b000000000000000000000110010000;
						 MAC7_W_I<=30'b111111111111111111100000100111;
						 MAC8_W_R<=0;
						 MAC8_W_I<=30'b111111111111111111100000000000;
						 MAC9_W_R<=30'b111111111111111111111001110000;
						 MAC9_W_I<=30'b111111111111111111100000100111;
						 MAC10_W_R<=30'b111111111111111111110011110000;
						 MAC10_W_I<=30'b111111111111111111100010011100;
						 MAC11_W_R<=30'b111111111111111111101110001110;
						 MAC11_W_I<=30'b111111111111111111100101011001;
						 MAC12_W_R<=30'b111111111111111111101001011000;
						 MAC12_W_I<=30'b111111111111111111101001011000;
						 MAC13_W_R<=30'b111111111111111111100101011001;
						 MAC13_W_I<=30'b111111111111111111101110001110;
						 MAC14_W_R<=30'b111111111111111111100010011100;
						 MAC14_W_I<=30'b111111111111111111110011110000;
						 MAC15_W_R<=30'b111111111111111111100000100111;
						 MAC15_W_I<=30'b111111111111111111111001110000;		
				end
			else 
				begin
						 MAC0_IN1_R<=0;
						 MAC0_IN1_I<=0;
						 MAC0_IN2_R<=0;
						 MAC0_IN2_I<=0;
						 MAC1_IN1_R<=0;
						 MAC1_IN1_I<=0;
						 MAC1_IN2_R<=0;
						 MAC1_IN2_I<=0;
						 MAC2_IN1_R<=0;
						 MAC2_IN1_I<=0;
						 MAC2_IN2_R<=0;
						 MAC2_IN2_I<=0;
						 MAC3_IN1_R<=0;
						 MAC3_IN1_I<=0;
						 MAC3_IN2_R<=0;
						 MAC3_IN2_I<=0;
						 MAC4_IN1_R<=0;
						 MAC4_IN1_I<=0;
						 MAC4_IN2_R<=0;
						 MAC4_IN2_I<=0;
						 MAC5_IN1_R<=0;
						 MAC5_IN1_I<=0;
						 MAC5_IN2_R<=0;
						 MAC5_IN2_I<=0;
						 MAC6_IN1_R<=0;
						 MAC6_IN1_I<=0;
						 MAC6_IN2_R<=0;
						 MAC6_IN2_I<=0;
						 MAC7_IN1_R<=0;
						 MAC7_IN1_I<=0;
						 MAC7_IN2_R<=0;
						 MAC7_IN2_I<=0;
						 MAC8_IN1_R<=0;
						 MAC8_IN1_I<=0;
						 MAC8_IN2_R<=0;
						 MAC8_IN2_I<=0;
						 MAC9_IN1_R<=0;
						 MAC9_IN1_I<=0;
						 MAC9_IN2_R<=0;
						 MAC9_IN2_I<=0;
						 MAC10_IN1_R<=0;
						 MAC10_IN1_I<=0;
						 MAC10_IN2_R<=0;
						 MAC10_IN2_I<=0;
						 MAC11_IN1_R<=0;
						 MAC11_IN1_I<=0;
						 MAC11_IN2_R<=0;
						 MAC11_IN2_I<=0;
						 MAC12_IN1_R<=0;
						 MAC12_IN1_I<=0;
						 MAC12_IN2_R<=0;
						 MAC12_IN2_I<=0;
						 MAC13_IN1_R<=0;
						 MAC13_IN1_I<=0;
						 MAC13_IN2_R<=0;
						 MAC13_IN2_I<=0;
						 MAC14_IN1_R<=0;
						 MAC14_IN1_I<=0;
						 MAC14_IN2_R<=0;
						 MAC14_IN2_I<=0;
						 MAC15_IN1_R<=0;
						 MAC15_IN1_I<=0;
						 MAC15_IN2_R<=0;
						 MAC15_IN2_I<=0;
						 
						 MAC0_W_R<=0;
						 MAC0_W_I<=0;
						 MAC1_W_R<=0;
						 MAC1_W_I<=0;
						 MAC2_W_R<=0;
						 MAC2_W_I<=0;
						 MAC3_W_R<=0;
						 MAC3_W_I<=0;
						 MAC4_W_R<=0;
						 MAC4_W_I<=0;
						 MAC5_W_R<=0;
						 MAC5_W_I<=0;
						 MAC6_W_R<=0;
						 MAC6_W_I<=0;
						 MAC7_W_R<=0;
						 MAC7_W_I<=0;
						 MAC8_W_R<=0;
						 MAC8_W_I<=0;
						 MAC9_W_R<=0;
						 MAC9_W_I<=0;
						 MAC10_W_R<=0;
						 MAC10_W_I<=0;
						 MAC11_W_R<=0;
						 MAC11_W_I<=0;
						 MAC12_W_R<=0;
						 MAC12_W_I<=0;
						 MAC13_W_R<=0;
						 MAC13_W_I<=0;
						 MAC14_W_R<=0;
						 MAC14_W_I<=0;
						 MAC15_W_R<=0;
						 MAC15_W_I<=0;	
				end
end
		
	
	
	
	// Control Unit 
	
	Control_Unit # () CU0
	(
		.CLK(CLK),
		.RST(RST),
		.EN(EN),
		.E0(E0),
		.E1(E1),
		.E2(E2),
		.E3(E3),
		.E4(E4),
		.S(Sel)
	);
	
	

	
	MAC # (.I(I) , .F(F)) MAC0
	(
		.IN1_R(MAC0_IN1_R),
		.IN1_I(MAC0_IN1_I),
		.IN2_R(MAC0_IN2_R),
		.IN2_I(MAC0_IN2_I),
		.W_R( MAC0_W_R),
		.W_I(MAC0_W_I),
		.OUT1_R(MAC0_OUT1_R),
		.OUT1_I(MAC0_OUT1_I),
		.OUT2_R(MAC0_OUT2_R),
		.OUT2_I(MAC0_OUT2_I)
	);
	
	
	MAC # (.I(I) , .F(F)) MAC1
	(
		.IN1_R(MAC1_IN1_R),
		.IN1_I(MAC1_IN1_I),
		.IN2_R(MAC1_IN2_R),
		.IN2_I(MAC1_IN2_I),
		.W_R( MAC1_W_R),
		.W_I(MAC1_W_I),
		.OUT1_R(MAC1_OUT1_R),
		.OUT1_I(MAC1_OUT1_I),
		.OUT2_R(MAC1_OUT2_R),
		.OUT2_I(MAC1_OUT2_I)
	);
	
	MAC # (.I(I) , .F(F)) MAC2
	(
		.IN1_R(MAC2_IN1_R),
		.IN1_I(MAC2_IN1_I),
		.IN2_R(MAC2_IN2_R),
		.IN2_I(MAC2_IN2_I),
		.W_R( MAC2_W_R),
		.W_I(MAC2_W_I),
		.OUT1_R(MAC2_OUT1_R),
		.OUT1_I(MAC2_OUT1_I),
		.OUT2_R(MAC2_OUT2_R),
		.OUT2_I(MAC2_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC3
	(
		.IN1_R(MAC3_IN1_R),
		.IN1_I(MAC3_IN1_I),
		.IN2_R(MAC3_IN2_R),
		.IN2_I(MAC3_IN2_I),
		.W_R( MAC3_W_R),
		.W_I(MAC3_W_I),
		.OUT1_R(MAC3_OUT1_R),
		.OUT1_I(MAC3_OUT1_I),
		.OUT2_R(MAC3_OUT2_R),
		.OUT2_I(MAC3_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC4
	(
		.IN1_R(MAC4_IN1_R),
		.IN1_I(MAC4_IN1_I),
		.IN2_R(MAC4_IN2_R),
		.IN2_I(MAC4_IN2_I),
		.W_R( MAC4_W_R),
		.W_I(MAC4_W_I),
		.OUT1_R(MAC4_OUT1_R),
		.OUT1_I(MAC4_OUT1_I),
		.OUT2_R(MAC4_OUT2_R),
		.OUT2_I(MAC4_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC5
	(
		.IN1_R(MAC5_IN1_R),
		.IN1_I(MAC5_IN1_I),
		.IN2_R(MAC5_IN2_R),
		.IN2_I(MAC5_IN2_I),
		.W_R( MAC5_W_R),
		.W_I(MAC5_W_I),
		.OUT1_R(MAC5_OUT1_R),
		.OUT1_I(MAC5_OUT1_I),
		.OUT2_R(MAC5_OUT2_R),
		.OUT2_I(MAC5_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC6
	(
		.IN1_R(MAC6_IN1_R),
		.IN1_I(MAC6_IN1_I),
		.IN2_R(MAC6_IN2_R),
		.IN2_I(MAC6_IN2_I),
		.W_R( MAC6_W_R),
		.W_I(MAC6_W_I),
		.OUT1_R(MAC6_OUT1_R),
		.OUT1_I(MAC6_OUT1_I),
		.OUT2_R(MAC6_OUT2_R),
		.OUT2_I(MAC6_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC7
	(
		.IN1_R(MAC7_IN1_R),
		.IN1_I(MAC7_IN1_I),
		.IN2_R(MAC7_IN2_R),
		.IN2_I(MAC7_IN2_I),
		.W_R( MAC7_W_R),
		.W_I(MAC7_W_I),
		.OUT1_R(MAC7_OUT1_R),
		.OUT1_I(MAC7_OUT1_I),
		.OUT2_R(MAC7_OUT2_R),
		.OUT2_I(MAC7_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC8
	(
		.IN1_R(MAC8_IN1_R),
		.IN1_I(MAC8_IN1_I),
		.IN2_R(MAC8_IN2_R),
		.IN2_I(MAC8_IN2_I),
		.W_R( MAC8_W_R),
		.W_I(MAC8_W_I),
		.OUT1_R(MAC8_OUT1_R),
		.OUT1_I(MAC8_OUT1_I),
		.OUT2_R(MAC8_OUT2_R),
		.OUT2_I(MAC8_OUT2_I)
	);
	
	MAC # (.I(I) , .F(F)) MAC9
	(
		.IN1_R(MAC9_IN1_R),
		.IN1_I(MAC9_IN1_I),
		.IN2_R(MAC9_IN2_R),
		.IN2_I(MAC9_IN2_I),
		.W_R( MAC9_W_R),
		.W_I(MAC9_W_I),
		.OUT1_R(MAC9_OUT1_R),
		.OUT1_I(MAC9_OUT1_I),
		.OUT2_R(MAC9_OUT2_R),
		.OUT2_I(MAC9_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC10
	(
		.IN1_R(MAC10_IN1_R),
		.IN1_I(MAC10_IN1_I),
		.IN2_R(MAC10_IN2_R),
		.IN2_I(MAC10_IN2_I),
		.W_R( MAC10_W_R),
		.W_I(MAC10_W_I),
		.OUT1_R(MAC10_OUT1_R),
		.OUT1_I(MAC10_OUT1_I),
		.OUT2_R(MAC10_OUT2_R),
		.OUT2_I(MAC10_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC11
	(
		.IN1_R(MAC11_IN1_R),
		.IN1_I(MAC11_IN1_I),
		.IN2_R(MAC11_IN2_R),
		.IN2_I(MAC11_IN2_I),
		.W_R( MAC11_W_R),
		.W_I(MAC11_W_I),
		.OUT1_R(MAC11_OUT1_R),
		.OUT1_I(MAC11_OUT1_I),
		.OUT2_R(MAC11_OUT2_R),
		.OUT2_I(MAC11_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC12
	(
		.IN1_R(MAC12_IN1_R),
		.IN1_I(MAC12_IN1_I),
		.IN2_R(MAC12_IN2_R),
		.IN2_I(MAC12_IN2_I),
		.W_R( MAC12_W_R),
		.W_I(MAC12_W_I),
		.OUT1_R(MAC12_OUT1_R),
		.OUT1_I(MAC12_OUT1_I),
		.OUT2_R(MAC12_OUT2_R),
		.OUT2_I(MAC12_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC13
	(
		.IN1_R(MAC13_IN1_R),
		.IN1_I(MAC13_IN1_I),
		.IN2_R(MAC13_IN2_R),
		.IN2_I(MAC13_IN2_I),
		.W_R( MAC13_W_R),
		.W_I(MAC13_W_I),
		.OUT1_R(MAC13_OUT1_R),
		.OUT1_I(MAC13_OUT1_I),
		.OUT2_R(MAC13_OUT2_R),
		.OUT2_I(MAC13_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC14
	(
		.IN1_R(MAC14_IN1_R),
		.IN1_I(MAC14_IN1_I),
		.IN2_R(MAC14_IN2_R),
		.IN2_I(MAC14_IN2_I),
		.W_R( MAC14_W_R),
		.W_I(MAC14_W_I),
		.OUT1_R(MAC14_OUT1_R),
		.OUT1_I(MAC14_OUT1_I),
		.OUT2_R(MAC14_OUT2_R),
		.OUT2_I(MAC14_OUT2_I)
	);

	MAC # (.I(I) , .F(F)) MAC15
	(
		.IN1_R(MAC15_IN1_R),
		.IN1_I(MAC15_IN1_I),
		.IN2_R(MAC15_IN2_R),
		.IN2_I(MAC15_IN2_I),
		.W_R( MAC15_W_R),
		.W_I(MAC15_W_I),
		.OUT1_R(MAC15_OUT1_R),
		.OUT1_I(MAC15_OUT1_I),
		.OUT2_R(MAC15_OUT2_R),
		.OUT2_I(MAC15_OUT2_I)
	);




	
	// Reg File
	
	Regfile# (.I(I) , .F(F)) RG0
	(
	.CLK (CLK),
	.RST (RST),
	.EN (E0),
	
	.IN_0_r (MAC0_OUT1_R),
	.IN_1_r (MAC0_OUT2_R),
	.IN_2_r (MAC1_OUT1_R),
	.IN_3_r (MAC1_OUT2_R),
	.IN_4_r (MAC2_OUT1_R),
	.IN_5_r (MAC2_OUT2_R),
	.IN_6_r (MAC3_OUT1_R),
	.IN_7_r (MAC3_OUT2_R),
	.IN_8_r (MAC4_OUT1_R),
	.IN_9_r (MAC4_OUT2_R),
	.IN_10_r (MAC5_OUT1_R),
	.IN_11_r (MAC5_OUT2_R),
	.IN_12_r (MAC6_OUT1_R),
	.IN_13_r (MAC6_OUT2_R),
	.IN_14_r (MAC7_OUT1_R),
	.IN_15_r (MAC7_OUT2_R),
	.IN_16_r (MAC8_OUT1_R),
	.IN_17_r (MAC8_OUT2_R),
	.IN_18_r (MAC9_OUT1_R),
	.IN_19_r (MAC9_OUT2_R),
	.IN_20_r (MAC10_OUT1_R),
	.IN_21_r (MAC10_OUT2_R),
	.IN_22_r (MAC11_OUT1_R),
	.IN_23_r (MAC11_OUT2_R),
	.IN_24_r (MAC12_OUT1_R),
	.IN_25_r (MAC12_OUT2_R),
	.IN_26_r (MAC13_OUT1_R),
	.IN_27_r (MAC13_OUT2_R),
	.IN_28_r (MAC14_OUT1_R),
	.IN_29_r (MAC14_OUT2_R),
	.IN_30_r (MAC15_OUT1_R),
	.IN_31_r (MAC15_OUT2_R),
	
	.IN_0_i (MAC0_OUT1_I),
	.IN_1_i (MAC0_OUT2_I),
	.IN_2_i (MAC1_OUT1_I),
	.IN_3_i (MAC1_OUT2_I),
	.IN_4_i (MAC2_OUT1_I),
	.IN_5_i (MAC2_OUT2_I),
	.IN_6_i (MAC3_OUT1_I),
	.IN_7_i (MAC3_OUT2_I),
	.IN_8_i (MAC4_OUT1_I),
	.IN_9_i (MAC4_OUT2_I),
	.IN_10_i (MAC5_OUT1_I),
	.IN_11_i (MAC5_OUT2_I),
	.IN_12_i (MAC6_OUT1_I),
	.IN_13_i (MAC6_OUT2_I),
	.IN_14_i (MAC7_OUT1_I),
	.IN_15_i (MAC7_OUT2_I),
	.IN_16_i (MAC8_OUT1_I),
	.IN_17_i (MAC8_OUT2_I),
	.IN_18_i (MAC9_OUT1_I),
	.IN_19_i (MAC9_OUT2_I),
	.IN_20_i (MAC10_OUT1_I),
	.IN_21_i (MAC10_OUT2_I),
	.IN_22_i (MAC11_OUT1_I),
	.IN_23_i (MAC11_OUT2_I),
	.IN_24_i (MAC12_OUT1_I),
	.IN_25_i (MAC12_OUT2_I),
	.IN_26_i (MAC13_OUT1_I),
	.IN_27_i (MAC13_OUT2_I),
	.IN_28_i (MAC14_OUT1_I),
	.IN_29_i (MAC14_OUT2_I),
	.IN_30_i (MAC15_OUT1_I),
	.IN_31_i (MAC15_OUT2_I),
	
	.OUT_0_r (regfile0_out0_r),
	.OUT_1_r (regfile0_out1_r),
	.OUT_2_r (regfile0_out2_r),
	.OUT_3_r (regfile0_out3_r),
	.OUT_4_r (regfile0_out4_r),
	.OUT_5_r (regfile0_out5_r),
	.OUT_6_r (regfile0_out6_r),
	.OUT_7_r (regfile0_out7_r),
	.OUT_8_r (regfile0_out8_r),
	.OUT_9_r (regfile0_out9_r),
	.OUT_10_r (regfile0_out10_r),
	.OUT_11_r (regfile0_out11_r),
	.OUT_12_r (regfile0_out12_r),
	.OUT_13_r (regfile0_out13_r),
	.OUT_14_r (regfile0_out14_r),
	.OUT_15_r (regfile0_out15_r),
	.OUT_16_r (regfile0_out16_r),
	.OUT_17_r (regfile0_out17_r),
	.OUT_18_r (regfile0_out18_r),
	.OUT_19_r (regfile0_out19_r),
	.OUT_20_r (regfile0_out20_r),
	.OUT_21_r (regfile0_out21_r),
	.OUT_22_r (regfile0_out22_r),
	.OUT_23_r (regfile0_out23_r),
	.OUT_24_r (regfile0_out24_r),
	.OUT_25_r (regfile0_out25_r),
	.OUT_26_r (regfile0_out26_r),
	.OUT_27_r (regfile0_out27_r),
	.OUT_28_r (regfile0_out28_r),
	.OUT_29_r (regfile0_out29_r),
	.OUT_30_r (regfile0_out30_r),
	.OUT_31_r (regfile0_out31_r),
	
	.OUT_0_i (regfile0_out0_i),
	.OUT_1_i (regfile0_out1_i),
	.OUT_2_i (regfile0_out2_i),
	.OUT_3_i (regfile0_out3_i),
	.OUT_4_i (regfile0_out4_i),
	.OUT_5_i (regfile0_out5_i),
	.OUT_6_i (regfile0_out6_i),
	.OUT_7_i (regfile0_out7_i),
	.OUT_8_i (regfile0_out8_i),
	.OUT_9_i (regfile0_out9_i),
	.OUT_10_i (regfile0_out10_i),
	.OUT_11_i (regfile0_out11_i),
	.OUT_12_i (regfile0_out12_i),
	.OUT_13_i (regfile0_out13_i),
	.OUT_14_i (regfile0_out14_i),
	.OUT_15_i (regfile0_out15_i),
	.OUT_16_i (regfile0_out16_i),
	.OUT_17_i (regfile0_out17_i),
	.OUT_18_i (regfile0_out18_i),
	.OUT_19_i (regfile0_out19_i),
	.OUT_20_i (regfile0_out20_i),
	.OUT_21_i (regfile0_out21_i),
	.OUT_22_i (regfile0_out22_i),
	.OUT_23_i (regfile0_out23_i),
	.OUT_24_i (regfile0_out24_i),
	.OUT_25_i (regfile0_out25_i),
	.OUT_26_i (regfile0_out26_i),
	.OUT_27_i (regfile0_out27_i),
	.OUT_28_i (regfile0_out28_i),
	.OUT_29_i (regfile0_out29_i),
	.OUT_30_i (regfile0_out30_i),
	.OUT_31_i (regfile0_out31_i)
	
	);
	



	Regfile # (.I(I) , .F(F)) RG1
	(
	.CLK (CLK),
	.RST (RST),
	.EN (E1),
	
	.IN_0_r (MAC0_OUT1_R),
	.IN_1_r (MAC1_OUT1_R),
	.IN_2_r (MAC0_OUT2_R),
	.IN_3_r (MAC1_OUT2_R),
	.IN_4_r (MAC2_OUT1_R),
	.IN_5_r (MAC3_OUT1_R),
	.IN_6_r (MAC2_OUT2_R),
	.IN_7_r (MAC3_OUT2_R),
	.IN_8_r (MAC4_OUT1_R),
	.IN_9_r (MAC5_OUT1_R),
	.IN_10_r (MAC4_OUT2_R),
	.IN_11_r (MAC5_OUT2_R),
	.IN_12_r (MAC6_OUT1_R),
	.IN_13_r (MAC7_OUT1_R),
	.IN_14_r (MAC6_OUT2_R),
	.IN_15_r (MAC7_OUT2_R),
	.IN_16_r (MAC8_OUT1_R),
	.IN_17_r (MAC9_OUT1_R),
	.IN_18_r (MAC8_OUT2_R),
	.IN_19_r (MAC9_OUT2_R),
	.IN_20_r (MAC10_OUT1_R),
	.IN_21_r (MAC11_OUT1_R),
	.IN_22_r (MAC10_OUT2_R),
	.IN_23_r (MAC11_OUT2_R),
	.IN_24_r (MAC12_OUT1_R),
	.IN_25_r (MAC13_OUT1_R),
	.IN_26_r (MAC12_OUT2_R),
	.IN_27_r (MAC13_OUT2_R),
	.IN_28_r (MAC14_OUT1_R),
	.IN_29_r (MAC15_OUT1_R),
	.IN_30_r (MAC14_OUT2_R),
	.IN_31_r (MAC15_OUT2_R),
	
	.IN_0_i (MAC0_OUT1_I),
	.IN_1_i (MAC1_OUT1_I),
	.IN_2_i (MAC0_OUT2_I),
	.IN_3_i (MAC1_OUT2_I),
	.IN_4_i (MAC2_OUT1_I),
	.IN_5_i (MAC3_OUT1_I),
	.IN_6_i (MAC2_OUT2_I),
	.IN_7_i (MAC3_OUT2_I),
	.IN_8_i (MAC4_OUT1_I),
	.IN_9_i (MAC5_OUT1_I),
	.IN_10_i (MAC4_OUT2_I),
	.IN_11_i (MAC5_OUT2_I),
	.IN_12_i (MAC6_OUT1_I),
	.IN_13_i (MAC7_OUT1_I),
	.IN_14_i (MAC6_OUT2_I),
	.IN_15_i (MAC7_OUT2_I),
	.IN_16_i (MAC8_OUT1_I),
	.IN_17_i (MAC9_OUT1_I),
	.IN_18_i (MAC8_OUT2_I),
	.IN_19_i (MAC9_OUT2_I),
	.IN_20_i (MAC10_OUT1_I),
	.IN_21_i (MAC11_OUT1_I),
	.IN_22_i (MAC10_OUT2_I),
	.IN_23_i (MAC11_OUT2_I),
	.IN_24_i (MAC12_OUT1_I),
	.IN_25_i (MAC13_OUT1_I),
	.IN_26_i (MAC12_OUT2_I),
	.IN_27_i (MAC13_OUT2_I),
	.IN_28_i (MAC14_OUT1_I),
	.IN_29_i (MAC15_OUT1_I),
	.IN_30_i (MAC14_OUT2_I),
	.IN_31_i (MAC15_OUT2_I),
	
	.OUT_0_r (regfile1_out0_r),
	.OUT_1_r (regfile1_out1_r),
	.OUT_2_r (regfile1_out2_r),
	.OUT_3_r (regfile1_out3_r),
	.OUT_4_r (regfile1_out4_r),
	.OUT_5_r (regfile1_out5_r),
	.OUT_6_r (regfile1_out6_r),
	.OUT_7_r (regfile1_out7_r),
	.OUT_8_r (regfile1_out8_r),
	.OUT_9_r (regfile1_out9_r),
	.OUT_10_r (regfile1_out10_r),
	.OUT_11_r (regfile1_out11_r),
	.OUT_12_r (regfile1_out12_r),
	.OUT_13_r (regfile1_out13_r),
	.OUT_14_r (regfile1_out14_r),
	.OUT_15_r (regfile1_out15_r),
	.OUT_16_r (regfile1_out16_r),
	.OUT_17_r (regfile1_out17_r),
	.OUT_18_r (regfile1_out18_r),
	.OUT_19_r (regfile1_out19_r),
	.OUT_20_r (regfile1_out20_r),
	.OUT_21_r (regfile1_out21_r),
	.OUT_22_r (regfile1_out22_r),
	.OUT_23_r (regfile1_out23_r),
	.OUT_24_r (regfile1_out24_r),
	.OUT_25_r (regfile1_out25_r),
	.OUT_26_r (regfile1_out26_r),
	.OUT_27_r (regfile1_out27_r),
	.OUT_28_r (regfile1_out28_r),
	.OUT_29_r (regfile1_out29_r),
	.OUT_30_r (regfile1_out30_r),
	.OUT_31_r (regfile1_out31_r),
	
	.OUT_0_i (regfile1_out0_i),
	.OUT_1_i (regfile1_out1_i),
	.OUT_2_i (regfile1_out2_i),
	.OUT_3_i (regfile1_out3_i),
	.OUT_4_i (regfile1_out4_i),
	.OUT_5_i (regfile1_out5_i),
	.OUT_6_i (regfile1_out6_i),
	.OUT_7_i (regfile1_out7_i),
	.OUT_8_i (regfile1_out8_i),
	.OUT_9_i (regfile1_out9_i),
	.OUT_10_i (regfile1_out10_i),
	.OUT_11_i (regfile1_out11_i),
	.OUT_12_i (regfile1_out12_i),
	.OUT_13_i (regfile1_out13_i),
	.OUT_14_i (regfile1_out14_i),
	.OUT_15_i (regfile1_out15_i),
	.OUT_16_i (regfile1_out16_i),
	.OUT_17_i (regfile1_out17_i),
	.OUT_18_i (regfile1_out18_i),
	.OUT_19_i (regfile1_out19_i),
	.OUT_20_i (regfile1_out20_i),
	.OUT_21_i (regfile1_out21_i),
	.OUT_22_i (regfile1_out22_i),
	.OUT_23_i (regfile1_out23_i),
	.OUT_24_i (regfile1_out24_i),
	.OUT_25_i (regfile1_out25_i),
	.OUT_26_i (regfile1_out26_i),
	.OUT_27_i (regfile1_out27_i),
	.OUT_28_i (regfile1_out28_i),
	.OUT_29_i (regfile1_out29_i),
	.OUT_30_i (regfile1_out30_i),
	.OUT_31_i (regfile1_out31_i)
	
	);
	
	
	
	
	Regfile # (.I(I) , .F(F)) RG2
	(
	.CLK (CLK),
	.RST (RST),
	.EN (E2),
	
	.IN_0_r (MAC0_OUT1_R),
	.IN_1_r (MAC1_OUT1_R),
	.IN_2_r (MAC2_OUT1_R),
	.IN_3_r (MAC3_OUT1_R),
	.IN_4_r (MAC0_OUT2_R),
	.IN_5_r (MAC1_OUT2_R),
	.IN_6_r (MAC2_OUT2_R),
	.IN_7_r (MAC3_OUT2_R),
	.IN_8_r (MAC4_OUT1_R),
	.IN_9_r (MAC5_OUT1_R),
	.IN_10_r (MAC6_OUT1_R),
	.IN_11_r (MAC7_OUT1_R),
	.IN_12_r (MAC4_OUT2_R),
	.IN_13_r (MAC5_OUT2_R),
	.IN_14_r (MAC6_OUT2_R),
	.IN_15_r (MAC7_OUT2_R),
	.IN_16_r (MAC8_OUT1_R),
	.IN_17_r (MAC9_OUT1_R),
	.IN_18_r (MAC10_OUT1_R),
	.IN_19_r (MAC11_OUT1_R),
	.IN_20_r (MAC8_OUT2_R),
	.IN_21_r (MAC9_OUT2_R),
	.IN_22_r (MAC10_OUT2_R),
	.IN_23_r (MAC11_OUT2_R),
	.IN_24_r (MAC12_OUT1_R),
	.IN_25_r (MAC13_OUT1_R),
	.IN_26_r (MAC14_OUT1_R),
	.IN_27_r (MAC15_OUT1_R),
	.IN_28_r (MAC12_OUT2_R),
	.IN_29_r (MAC13_OUT2_R),
	.IN_30_r (MAC14_OUT2_R),
	.IN_31_r (MAC15_OUT2_R),
	
	.IN_0_i (MAC0_OUT1_I),
	.IN_1_i (MAC1_OUT1_I),
	.IN_2_i (MAC2_OUT1_I),
	.IN_3_i (MAC3_OUT1_I),
	.IN_4_i (MAC0_OUT2_I),
	.IN_5_i (MAC1_OUT2_I),
	.IN_6_i (MAC2_OUT2_I),
	.IN_7_i (MAC3_OUT2_I),
	.IN_8_i (MAC4_OUT1_I),
	.IN_9_i (MAC5_OUT1_I),
	.IN_10_i (MAC6_OUT1_I),
	.IN_11_i (MAC7_OUT1_I),
	.IN_12_i (MAC4_OUT2_I),
	.IN_13_i (MAC5_OUT2_I),
	.IN_14_i (MAC6_OUT2_I),
	.IN_15_i (MAC7_OUT2_I),
	.IN_16_i (MAC8_OUT1_I),
	.IN_17_i (MAC9_OUT1_I),
	.IN_18_i (MAC10_OUT1_I),
	.IN_19_i (MAC11_OUT1_I),
	.IN_20_i (MAC8_OUT2_I),
	.IN_21_i (MAC9_OUT2_I),
	.IN_22_i (MAC10_OUT2_I),
	.IN_23_i (MAC11_OUT2_I),
	.IN_24_i (MAC12_OUT1_I),
	.IN_25_i (MAC13_OUT1_I),
	.IN_26_i (MAC14_OUT1_I),
	.IN_27_i (MAC15_OUT1_I),
	.IN_28_i (MAC12_OUT2_I),
	.IN_29_i (MAC13_OUT2_I),
	.IN_30_i (MAC14_OUT2_I),
	.IN_31_i (MAC15_OUT2_I),
	
	.OUT_0_r (regfile2_out0_r),
	.OUT_1_r (regfile2_out1_r),
	.OUT_2_r (regfile2_out2_r),
	.OUT_3_r (regfile2_out3_r),
	.OUT_4_r (regfile2_out4_r),
	.OUT_5_r (regfile2_out5_r),
	.OUT_6_r (regfile2_out6_r),
	.OUT_7_r (regfile2_out7_r),
	.OUT_8_r (regfile2_out8_r),
	.OUT_9_r (regfile2_out9_r),
	.OUT_10_r (regfile2_out10_r),
	.OUT_11_r (regfile2_out11_r),
	.OUT_12_r (regfile2_out12_r),
	.OUT_13_r (regfile2_out13_r),
	.OUT_14_r (regfile2_out14_r),
	.OUT_15_r (regfile2_out15_r),
	.OUT_16_r (regfile2_out16_r),
	.OUT_17_r (regfile2_out17_r),
	.OUT_18_r (regfile2_out18_r),
	.OUT_19_r (regfile2_out19_r),
	.OUT_20_r (regfile2_out20_r),
	.OUT_21_r (regfile2_out21_r),
	.OUT_22_r (regfile2_out22_r),
	.OUT_23_r (regfile2_out23_r),
	.OUT_24_r (regfile2_out24_r),
	.OUT_25_r (regfile2_out25_r),
	.OUT_26_r (regfile2_out26_r),
	.OUT_27_r (regfile2_out27_r),
	.OUT_28_r (regfile2_out28_r),
	.OUT_29_r (regfile2_out29_r),
	.OUT_30_r (regfile2_out30_r),
	.OUT_31_r (regfile2_out31_r),
	
	.OUT_0_i (regfile2_out0_i),
	.OUT_1_i (regfile2_out1_i),
	.OUT_2_i (regfile2_out2_i),
	.OUT_3_i (regfile2_out3_i),
	.OUT_4_i (regfile2_out4_i),
	.OUT_5_i (regfile2_out5_i),
	.OUT_6_i (regfile2_out6_i),
	.OUT_7_i (regfile2_out7_i),
	.OUT_8_i (regfile2_out8_i),
	.OUT_9_i (regfile2_out9_i),
	.OUT_10_i (regfile2_out10_i),
	.OUT_11_i (regfile2_out11_i),
	.OUT_12_i (regfile2_out12_i),
	.OUT_13_i (regfile2_out13_i),
	.OUT_14_i (regfile2_out14_i),
	.OUT_15_i (regfile2_out15_i),
	.OUT_16_i (regfile2_out16_i),
	.OUT_17_i (regfile2_out17_i),
	.OUT_18_i (regfile2_out18_i),
	.OUT_19_i (regfile2_out19_i),
	.OUT_20_i (regfile2_out20_i),
	.OUT_21_i (regfile2_out21_i),
	.OUT_22_i (regfile2_out22_i),
	.OUT_23_i (regfile2_out23_i),
	.OUT_24_i (regfile2_out24_i),
	.OUT_25_i (regfile2_out25_i),
	.OUT_26_i (regfile2_out26_i),
	.OUT_27_i (regfile2_out27_i),
	.OUT_28_i (regfile2_out28_i),
	.OUT_29_i (regfile2_out29_i),
	.OUT_30_i (regfile2_out30_i),
	.OUT_31_i (regfile2_out31_i)
	
	);
	
	
	
	Regfile # (.I(I) , .F(F)) RG3
	(
	.CLK (CLK),
	.RST (RST),
	.EN (E3),
	.IN_0_r (MAC0_OUT1_R),
	.IN_1_r (MAC1_OUT1_R),
	.IN_2_r (MAC2_OUT1_R),
	.IN_3_r (MAC3_OUT1_R),
	.IN_4_r (MAC4_OUT1_R),
	.IN_5_r (MAC5_OUT1_R),
	.IN_6_r (MAC6_OUT1_R),
	.IN_7_r (MAC7_OUT1_R),
	.IN_8_r (MAC0_OUT2_R),
	.IN_9_r (MAC1_OUT2_R),
	.IN_10_r (MAC2_OUT2_R),
	.IN_11_r (MAC3_OUT2_R),
	.IN_12_r (MAC4_OUT2_R),
	.IN_13_r (MAC5_OUT2_R),
	.IN_14_r (MAC6_OUT2_R),
	.IN_15_r (MAC7_OUT2_R),
	.IN_16_r (MAC8_OUT1_R),
	.IN_17_r (MAC9_OUT1_R),
	.IN_18_r (MAC10_OUT1_R),
	.IN_19_r (MAC11_OUT1_R),
	.IN_20_r (MAC12_OUT1_R),
	.IN_21_r (MAC13_OUT1_R),
	.IN_22_r (MAC14_OUT1_R),
	.IN_23_r (MAC15_OUT1_R),
	.IN_24_r (MAC8_OUT2_R),
	.IN_25_r (MAC9_OUT2_R),
	.IN_26_r (MAC10_OUT2_R),
	.IN_27_r (MAC11_OUT2_R),
	.IN_28_r (MAC12_OUT2_R),
	.IN_29_r (MAC13_OUT2_R),
	.IN_30_r (MAC14_OUT2_R),
	.IN_31_r (MAC15_OUT2_R),
	
	.IN_0_i (MAC0_OUT1_I),
	.IN_1_i (MAC1_OUT1_I),
	.IN_2_i (MAC2_OUT1_I),
	.IN_3_i (MAC3_OUT1_I),
	.IN_4_i (MAC4_OUT1_I),
	.IN_5_i (MAC5_OUT1_I),
	.IN_6_i (MAC6_OUT1_I),
	.IN_7_i (MAC7_OUT1_I),
	.IN_8_i (MAC0_OUT2_I),
	.IN_9_i (MAC1_OUT2_I),
	.IN_10_i (MAC2_OUT2_I),
	.IN_11_i (MAC3_OUT2_I),
	.IN_12_i (MAC4_OUT2_I),
	.IN_13_i (MAC5_OUT2_I),
	.IN_14_i (MAC6_OUT2_I),
	.IN_15_i (MAC7_OUT2_I),
	.IN_16_i (MAC8_OUT1_I),
	.IN_17_i (MAC9_OUT1_I),
	.IN_18_i (MAC10_OUT1_I),
	.IN_19_i (MAC11_OUT1_I),
	.IN_20_i (MAC12_OUT1_I),
	.IN_21_i (MAC13_OUT1_I),
	.IN_22_i (MAC14_OUT1_I),
	.IN_23_i (MAC15_OUT1_I),
	.IN_24_i (MAC8_OUT2_I),
	.IN_25_i (MAC9_OUT2_I),
	.IN_26_i (MAC10_OUT2_I),
	.IN_27_i (MAC11_OUT2_I),
	.IN_28_i (MAC12_OUT2_I),
	.IN_29_i (MAC13_OUT2_I),
	.IN_30_i (MAC14_OUT2_I),
	.IN_31_i (MAC15_OUT2_I),
	
	
	.OUT_0_r (regfile3_out0_r),
	.OUT_1_r (regfile3_out1_r),
	.OUT_2_r (regfile3_out2_r),
	.OUT_3_r (regfile3_out3_r),
	.OUT_4_r (regfile3_out4_r),
	.OUT_5_r (regfile3_out5_r),
	.OUT_6_r (regfile3_out6_r),
	.OUT_7_r (regfile3_out7_r),
	.OUT_8_r (regfile3_out8_r),
	.OUT_9_r (regfile3_out9_r),
	.OUT_10_r (regfile3_out10_r),
	.OUT_11_r (regfile3_out11_r),
	.OUT_12_r (regfile3_out12_r),
	.OUT_13_r (regfile3_out13_r),
	.OUT_14_r (regfile3_out14_r),
	.OUT_15_r (regfile3_out15_r),
	.OUT_16_r (regfile3_out16_r),
	.OUT_17_r (regfile3_out17_r),
	.OUT_18_r (regfile3_out18_r),
	.OUT_19_r (regfile3_out19_r),
	.OUT_20_r (regfile3_out20_r),
	.OUT_21_r (regfile3_out21_r),
	.OUT_22_r (regfile3_out22_r),
	.OUT_23_r (regfile3_out23_r),
	.OUT_24_r (regfile3_out24_r),
	.OUT_25_r (regfile3_out25_r),
	.OUT_26_r (regfile3_out26_r),
	.OUT_27_r (regfile3_out27_r),
	.OUT_28_r (regfile3_out28_r),
	.OUT_29_r (regfile3_out29_r),
	.OUT_30_r (regfile3_out30_r),
	.OUT_31_r (regfile3_out31_r),
	
	.OUT_0_i (regfile3_out0_i),
	.OUT_1_i (regfile3_out1_i),
	.OUT_2_i (regfile3_out2_i),
	.OUT_3_i (regfile3_out3_i),
	.OUT_4_i (regfile3_out4_i),
	.OUT_5_i (regfile3_out5_i),
	.OUT_6_i (regfile3_out6_i),
	.OUT_7_i (regfile3_out7_i),
	.OUT_8_i (regfile3_out8_i),
	.OUT_9_i (regfile3_out9_i),
	.OUT_10_i (regfile3_out10_i),
	.OUT_11_i (regfile3_out11_i),
	.OUT_12_i (regfile3_out12_i),
	.OUT_13_i (regfile3_out13_i),
	.OUT_14_i (regfile3_out14_i),
	.OUT_15_i (regfile3_out15_i),
	.OUT_16_i (regfile3_out16_i),
	.OUT_17_i (regfile3_out17_i),
	.OUT_18_i (regfile3_out18_i),
	.OUT_19_i (regfile3_out19_i),
	.OUT_20_i (regfile3_out20_i),
	.OUT_21_i (regfile3_out21_i),
	.OUT_22_i (regfile3_out22_i),
	.OUT_23_i (regfile3_out23_i),
	.OUT_24_i (regfile3_out24_i),
	.OUT_25_i (regfile3_out25_i),
	.OUT_26_i (regfile3_out26_i),
	.OUT_27_i (regfile3_out27_i),
	.OUT_28_i (regfile3_out28_i),
	.OUT_29_i (regfile3_out29_i),
	.OUT_30_i (regfile3_out30_i),
	.OUT_31_i (regfile3_out31_i)
	
	);
	
	
	
	Regfile # (.I(I) , .F(F)) RG4
	(
	.CLK (CLK),
	.RST (RST),
	.EN (E4),
	.IN_0_r (MAC0_OUT1_R),
	.IN_1_r (MAC0_OUT2_R),
	.IN_2_r (MAC1_OUT1_R),
	.IN_3_r (MAC1_OUT2_R),
	.IN_4_r (MAC2_OUT1_R),
	.IN_5_r (MAC2_OUT2_R),
	.IN_6_r (MAC3_OUT2_R),
	.IN_7_r (MAC3_OUT1_R),
	.IN_8_r (MAC4_OUT1_R),
	.IN_9_r (MAC4_OUT2_R),
	.IN_10_r (MAC5_OUT1_R),
	.IN_11_r (MAC5_OUT2_R),
	.IN_12_r (MAC6_OUT1_R),
	.IN_13_r (MAC6_OUT2_R),
	.IN_14_r (MAC7_OUT1_R),
	.IN_15_r (MAC7_OUT2_R),
	.IN_16_r (MAC8_OUT1_R),
	.IN_17_r (MAC8_OUT2_R),
	.IN_18_r (MAC9_OUT1_R),
	.IN_19_r (MAC9_OUT2_R),
	.IN_20_r (MAC10_OUT1_R),
	.IN_21_r (MAC10_OUT2_R),
	.IN_22_r (MAC11_OUT1_R),
	.IN_23_r (MAC11_OUT2_R),
	.IN_24_r (MAC12_OUT1_R),
	.IN_25_r (MAC12_OUT2_R),
	.IN_26_r (MAC13_OUT1_R),
	.IN_27_r (MAC13_OUT2_R),
	.IN_28_r (MAC14_OUT1_R),
	.IN_29_r (MAC14_OUT2_R),
	.IN_30_r (MAC15_OUT1_R),
	.IN_31_r (MAC15_OUT2_R),
	
	.IN_0_i (MAC0_OUT1_I),
	.IN_1_i (MAC0_OUT2_I),
	.IN_2_i (MAC1_OUT1_I),
	.IN_3_i (MAC1_OUT2_I),
	.IN_4_i (MAC2_OUT1_I),
	.IN_5_i (MAC2_OUT2_I),
	.IN_6_i (MAC3_OUT2_I),
	.IN_7_i (MAC3_OUT1_I),
	.IN_8_i (MAC4_OUT1_I),
	.IN_9_i (MAC4_OUT2_I),
	.IN_10_i (MAC5_OUT1_I),
	.IN_11_i (MAC5_OUT2_I),
	.IN_12_i (MAC6_OUT1_I),
	.IN_13_i (MAC6_OUT2_I),
	.IN_14_i (MAC7_OUT1_I),
	.IN_15_i (MAC7_OUT2_I),
	.IN_16_i (MAC8_OUT1_I),
	.IN_17_i (MAC8_OUT2_I),
	.IN_18_i (MAC9_OUT1_I),
	.IN_19_i (MAC9_OUT2_I),
	.IN_20_i (MAC10_OUT1_I),
	.IN_21_i (MAC10_OUT2_I),
	.IN_22_i (MAC11_OUT1_I),
	.IN_23_i (MAC11_OUT2_I),
	.IN_24_i (MAC12_OUT1_I),
	.IN_25_i (MAC12_OUT2_I),
	.IN_26_i (MAC13_OUT1_I),
	.IN_27_i (MAC13_OUT2_I),
	.IN_28_i (MAC14_OUT1_I),
	.IN_29_i (MAC14_OUT2_I),
	.IN_30_i (MAC15_OUT1_I),
	.IN_31_i (MAC15_OUT2_I),
	
	
	.OUT_0_r (OUT0_r),
	.OUT_1_r (OUT1_r),
	.OUT_2_r (OUT2_r),
	.OUT_3_r (OUT3_r),
	.OUT_4_r (OUT4_r),
	.OUT_5_r (OUT5_r),
	.OUT_6_r (OUT6_r),
	.OUT_7_r (OUT7_r),
	.OUT_8_r (OUT8_r),
	.OUT_9_r (OUT9_r),
	.OUT_10_r (OUT10_r),
	.OUT_11_r (OUT11_r),
	.OUT_12_r (OUT12_r),
	.OUT_13_r (OUT13_r),
	.OUT_14_r (OUT14_r),
	.OUT_15_r (OUT15_r),
	.OUT_16_r (OUT16_r),
	.OUT_17_r (OUT17_r),
	.OUT_18_r (OUT18_r),
	.OUT_19_r (OUT19_r),
	.OUT_20_r (OUT20_r),
	.OUT_21_r (OUT21_r),
	.OUT_22_r (OUT22_r),
	.OUT_23_r (OUT23_r),
	.OUT_24_r (OUT24_r),
	.OUT_25_r (OUT25_r),
	.OUT_26_r (OUT26_r),
	.OUT_27_r (OUT27_r),
	.OUT_28_r (OUT28_r),
	.OUT_29_r (OUT29_r),
	.OUT_30_r (OUT30_r),
	.OUT_31_r (OUT31_r),
	
	.OUT_0_i (OUT0_i),
	.OUT_1_i (OUT1_i),
	.OUT_2_i (OUT2_i),
	.OUT_3_i (OUT3_i),
	.OUT_4_i (OUT4_i),
	.OUT_5_i (OUT5_i),
	.OUT_6_i (OUT6_i),
	.OUT_7_i (OUT7_i),
	.OUT_8_i (OUT8_i),
	.OUT_9_i (OUT9_i),
	.OUT_10_i (OUT10_i),
	.OUT_11_i (OUT11_i),
	.OUT_12_i (OUT12_i),
	.OUT_13_i (OUT13_i),
	.OUT_14_i (OUT14_i),
	.OUT_15_i (OUT15_i),
	.OUT_16_i (OUT16_i),
	.OUT_17_i (OUT17_i),
	.OUT_18_i (OUT18_i),
	.OUT_19_i (OUT19_i),
	.OUT_20_i (OUT20_i),
	.OUT_21_i (OUT21_i),
	.OUT_22_i (OUT22_i),
	.OUT_23_i (OUT23_i),
	.OUT_24_i (OUT24_i),
	.OUT_25_i (OUT25_i),
	.OUT_26_i (OUT26_i),
	.OUT_27_i (OUT27_i),
	.OUT_28_i (OUT28_i),
	.OUT_29_i (OUT29_i),
	.OUT_30_i (OUT30_i),
	.OUT_31_i(OUT31_i)
	
	);
	
	
endmodule 